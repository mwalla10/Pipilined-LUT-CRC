module crctab_ev17
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h8167d675 ;
    mem[8'h2] <= 32'h60eb15d ;
    mem[8'h3] <= 32'h87696728 ;
    mem[8'h4] <= 32'hc1d62ba ;
    mem[8'h5] <= 32'h8d7ab4cf ;
    mem[8'h6] <= 32'ha13d3e7 ;
    mem[8'h7] <= 32'h8b740592 ;
    mem[8'h8] <= 32'h183ac574 ;
    mem[8'h9] <= 32'h995d1301 ;
    mem[8'ha] <= 32'h1e347429 ;
    mem[8'hb] <= 32'h9f53a25c ;
    mem[8'hc] <= 32'h1427a7ce ;
    mem[8'hd] <= 32'h954071bb ;
    mem[8'he] <= 32'h12291693 ;
    mem[8'hf] <= 32'h934ec0e6 ;
    mem[8'h10] <= 32'h30758ae8 ;
    mem[8'h11] <= 32'hb1125c9d ;
    mem[8'h12] <= 32'h367b3bb5 ;
    mem[8'h13] <= 32'hb71cedc0 ;
    mem[8'h14] <= 32'h3c68e852 ;
    mem[8'h15] <= 32'hbd0f3e27 ;
    mem[8'h16] <= 32'h3a66590f ;
    mem[8'h17] <= 32'hbb018f7a ;
    mem[8'h18] <= 32'h284f4f9c ;
    mem[8'h19] <= 32'ha92899e9 ;
    mem[8'h1a] <= 32'h2e41fec1 ;
    mem[8'h1b] <= 32'haf2628b4 ;
    mem[8'h1c] <= 32'h24522d26 ;
    mem[8'h1d] <= 32'ha535fb53 ;
    mem[8'h1e] <= 32'h225c9c7b ;
    mem[8'h1f] <= 32'ha33b4a0e ;
    mem[8'h20] <= 32'h60eb15d0 ;
    mem[8'h21] <= 32'he18cc3a5 ;
    mem[8'h22] <= 32'h66e5a48d ;
    mem[8'h23] <= 32'he78272f8 ;
    mem[8'h24] <= 32'h6cf6776a ;
    mem[8'h25] <= 32'hed91a11f ;
    mem[8'h26] <= 32'h6af8c637 ;
    mem[8'h27] <= 32'heb9f1042 ;
    mem[8'h28] <= 32'h78d1d0a4 ;
    mem[8'h29] <= 32'hf9b606d1 ;
    mem[8'h2a] <= 32'h7edf61f9 ;
    mem[8'h2b] <= 32'hffb8b78c ;
    mem[8'h2c] <= 32'h74ccb21e ;
    mem[8'h2d] <= 32'hf5ab646b ;
    mem[8'h2e] <= 32'h72c20343 ;
    mem[8'h2f] <= 32'hf3a5d536 ;
    mem[8'h30] <= 32'h509e9f38 ;
    mem[8'h31] <= 32'hd1f9494d ;
    mem[8'h32] <= 32'h56902e65 ;
    mem[8'h33] <= 32'hd7f7f810 ;
    mem[8'h34] <= 32'h5c83fd82 ;
    mem[8'h35] <= 32'hdde42bf7 ;
    mem[8'h36] <= 32'h5a8d4cdf ;
    mem[8'h37] <= 32'hdbea9aaa ;
    mem[8'h38] <= 32'h48a45a4c ;
    mem[8'h39] <= 32'hc9c38c39 ;
    mem[8'h3a] <= 32'h4eaaeb11 ;
    mem[8'h3b] <= 32'hcfcd3d64 ;
    mem[8'h3c] <= 32'h44b938f6 ;
    mem[8'h3d] <= 32'hc5deee83 ;
    mem[8'h3e] <= 32'h42b789ab ;
    mem[8'h3f] <= 32'hc3d05fde ;
    mem[8'h40] <= 32'hc1d62ba0 ;
    mem[8'h41] <= 32'h40b1fdd5 ;
    mem[8'h42] <= 32'hc7d89afd ;
    mem[8'h43] <= 32'h46bf4c88 ;
    mem[8'h44] <= 32'hcdcb491a ;
    mem[8'h45] <= 32'h4cac9f6f ;
    mem[8'h46] <= 32'hcbc5f847 ;
    mem[8'h47] <= 32'h4aa22e32 ;
    mem[8'h48] <= 32'hd9eceed4 ;
    mem[8'h49] <= 32'h588b38a1 ;
    mem[8'h4a] <= 32'hdfe25f89 ;
    mem[8'h4b] <= 32'h5e8589fc ;
    mem[8'h4c] <= 32'hd5f18c6e ;
    mem[8'h4d] <= 32'h54965a1b ;
    mem[8'h4e] <= 32'hd3ff3d33 ;
    mem[8'h4f] <= 32'h5298eb46 ;
    mem[8'h50] <= 32'hf1a3a148 ;
    mem[8'h51] <= 32'h70c4773d ;
    mem[8'h52] <= 32'hf7ad1015 ;
    mem[8'h53] <= 32'h76cac660 ;
    mem[8'h54] <= 32'hfdbec3f2 ;
    mem[8'h55] <= 32'h7cd91587 ;
    mem[8'h56] <= 32'hfbb072af ;
    mem[8'h57] <= 32'h7ad7a4da ;
    mem[8'h58] <= 32'he999643c ;
    mem[8'h59] <= 32'h68feb249 ;
    mem[8'h5a] <= 32'hef97d561 ;
    mem[8'h5b] <= 32'h6ef00314 ;
    mem[8'h5c] <= 32'he5840686 ;
    mem[8'h5d] <= 32'h64e3d0f3 ;
    mem[8'h5e] <= 32'he38ab7db ;
    mem[8'h5f] <= 32'h62ed61ae ;
    mem[8'h60] <= 32'ha13d3e70 ;
    mem[8'h61] <= 32'h205ae805 ;
    mem[8'h62] <= 32'ha7338f2d ;
    mem[8'h63] <= 32'h26545958 ;
    mem[8'h64] <= 32'had205cca ;
    mem[8'h65] <= 32'h2c478abf ;
    mem[8'h66] <= 32'hab2eed97 ;
    mem[8'h67] <= 32'h2a493be2 ;
    mem[8'h68] <= 32'hb907fb04 ;
    mem[8'h69] <= 32'h38602d71 ;
    mem[8'h6a] <= 32'hbf094a59 ;
    mem[8'h6b] <= 32'h3e6e9c2c ;
    mem[8'h6c] <= 32'hb51a99be ;
    mem[8'h6d] <= 32'h347d4fcb ;
    mem[8'h6e] <= 32'hb31428e3 ;
    mem[8'h6f] <= 32'h3273fe96 ;
    mem[8'h70] <= 32'h9148b498 ;
    mem[8'h71] <= 32'h102f62ed ;
    mem[8'h72] <= 32'h974605c5 ;
    mem[8'h73] <= 32'h1621d3b0 ;
    mem[8'h74] <= 32'h9d55d622 ;
    mem[8'h75] <= 32'h1c320057 ;
    mem[8'h76] <= 32'h9b5b677f ;
    mem[8'h77] <= 32'h1a3cb10a ;
    mem[8'h78] <= 32'h897271ec ;
    mem[8'h79] <= 32'h815a799 ;
    mem[8'h7a] <= 32'h8f7cc0b1 ;
    mem[8'h7b] <= 32'he1b16c4 ;
    mem[8'h7c] <= 32'h856f1356 ;
    mem[8'h7d] <= 32'h408c523 ;
    mem[8'h7e] <= 32'h8361a20b ;
    mem[8'h7f] <= 32'h206747e ;
    mem[8'h80] <= 32'h876d4af7 ;
    mem[8'h81] <= 32'h60a9c82 ;
    mem[8'h82] <= 32'h8163fbaa ;
    mem[8'h83] <= 32'h42ddf ;
    mem[8'h84] <= 32'h8b70284d ;
    mem[8'h85] <= 32'ha17fe38 ;
    mem[8'h86] <= 32'h8d7e9910 ;
    mem[8'h87] <= 32'hc194f65 ;
    mem[8'h88] <= 32'h9f578f83 ;
    mem[8'h89] <= 32'h1e3059f6 ;
    mem[8'h8a] <= 32'h99593ede ;
    mem[8'h8b] <= 32'h183ee8ab ;
    mem[8'h8c] <= 32'h934aed39 ;
    mem[8'h8d] <= 32'h122d3b4c ;
    mem[8'h8e] <= 32'h95445c64 ;
    mem[8'h8f] <= 32'h14238a11 ;
    mem[8'h90] <= 32'hb718c01f ;
    mem[8'h91] <= 32'h367f166a ;
    mem[8'h92] <= 32'hb1167142 ;
    mem[8'h93] <= 32'h3071a737 ;
    mem[8'h94] <= 32'hbb05a2a5 ;
    mem[8'h95] <= 32'h3a6274d0 ;
    mem[8'h96] <= 32'hbd0b13f8 ;
    mem[8'h97] <= 32'h3c6cc58d ;
    mem[8'h98] <= 32'haf22056b ;
    mem[8'h99] <= 32'h2e45d31e ;
    mem[8'h9a] <= 32'ha92cb436 ;
    mem[8'h9b] <= 32'h284b6243 ;
    mem[8'h9c] <= 32'ha33f67d1 ;
    mem[8'h9d] <= 32'h2258b1a4 ;
    mem[8'h9e] <= 32'ha531d68c ;
    mem[8'h9f] <= 32'h245600f9 ;
    mem[8'ha0] <= 32'he7865f27 ;
    mem[8'ha1] <= 32'h66e18952 ;
    mem[8'ha2] <= 32'he188ee7a ;
    mem[8'ha3] <= 32'h60ef380f ;
    mem[8'ha4] <= 32'heb9b3d9d ;
    mem[8'ha5] <= 32'h6afcebe8 ;
    mem[8'ha6] <= 32'hed958cc0 ;
    mem[8'ha7] <= 32'h6cf25ab5 ;
    mem[8'ha8] <= 32'hffbc9a53 ;
    mem[8'ha9] <= 32'h7edb4c26 ;
    mem[8'haa] <= 32'hf9b22b0e ;
    mem[8'hab] <= 32'h78d5fd7b ;
    mem[8'hac] <= 32'hf3a1f8e9 ;
    mem[8'had] <= 32'h72c62e9c ;
    mem[8'hae] <= 32'hf5af49b4 ;
    mem[8'haf] <= 32'h74c89fc1 ;
    mem[8'hb0] <= 32'hd7f3d5cf ;
    mem[8'hb1] <= 32'h569403ba ;
    mem[8'hb2] <= 32'hd1fd6492 ;
    mem[8'hb3] <= 32'h509ab2e7 ;
    mem[8'hb4] <= 32'hdbeeb775 ;
    mem[8'hb5] <= 32'h5a896100 ;
    mem[8'hb6] <= 32'hdde00628 ;
    mem[8'hb7] <= 32'h5c87d05d ;
    mem[8'hb8] <= 32'hcfc910bb ;
    mem[8'hb9] <= 32'h4eaec6ce ;
    mem[8'hba] <= 32'hc9c7a1e6 ;
    mem[8'hbb] <= 32'h48a07793 ;
    mem[8'hbc] <= 32'hc3d47201 ;
    mem[8'hbd] <= 32'h42b3a474 ;
    mem[8'hbe] <= 32'hc5dac35c ;
    mem[8'hbf] <= 32'h44bd1529 ;
    mem[8'hc0] <= 32'h46bb6157 ;
    mem[8'hc1] <= 32'hc7dcb722 ;
    mem[8'hc2] <= 32'h40b5d00a ;
    mem[8'hc3] <= 32'hc1d2067f ;
    mem[8'hc4] <= 32'h4aa603ed ;
    mem[8'hc5] <= 32'hcbc1d598 ;
    mem[8'hc6] <= 32'h4ca8b2b0 ;
    mem[8'hc7] <= 32'hcdcf64c5 ;
    mem[8'hc8] <= 32'h5e81a423 ;
    mem[8'hc9] <= 32'hdfe67256 ;
    mem[8'hca] <= 32'h588f157e ;
    mem[8'hcb] <= 32'hd9e8c30b ;
    mem[8'hcc] <= 32'h529cc699 ;
    mem[8'hcd] <= 32'hd3fb10ec ;
    mem[8'hce] <= 32'h549277c4 ;
    mem[8'hcf] <= 32'hd5f5a1b1 ;
    mem[8'hd0] <= 32'h76ceebbf ;
    mem[8'hd1] <= 32'hf7a93dca ;
    mem[8'hd2] <= 32'h70c05ae2 ;
    mem[8'hd3] <= 32'hf1a78c97 ;
    mem[8'hd4] <= 32'h7ad38905 ;
    mem[8'hd5] <= 32'hfbb45f70 ;
    mem[8'hd6] <= 32'h7cdd3858 ;
    mem[8'hd7] <= 32'hfdbaee2d ;
    mem[8'hd8] <= 32'h6ef42ecb ;
    mem[8'hd9] <= 32'hef93f8be ;
    mem[8'hda] <= 32'h68fa9f96 ;
    mem[8'hdb] <= 32'he99d49e3 ;
    mem[8'hdc] <= 32'h62e94c71 ;
    mem[8'hdd] <= 32'he38e9a04 ;
    mem[8'hde] <= 32'h64e7fd2c ;
    mem[8'hdf] <= 32'he5802b59 ;
    mem[8'he0] <= 32'h26507487 ;
    mem[8'he1] <= 32'ha737a2f2 ;
    mem[8'he2] <= 32'h205ec5da ;
    mem[8'he3] <= 32'ha13913af ;
    mem[8'he4] <= 32'h2a4d163d ;
    mem[8'he5] <= 32'hab2ac048 ;
    mem[8'he6] <= 32'h2c43a760 ;
    mem[8'he7] <= 32'had247115 ;
    mem[8'he8] <= 32'h3e6ab1f3 ;
    mem[8'he9] <= 32'hbf0d6786 ;
    mem[8'hea] <= 32'h386400ae ;
    mem[8'heb] <= 32'hb903d6db ;
    mem[8'hec] <= 32'h3277d349 ;
    mem[8'hed] <= 32'hb310053c ;
    mem[8'hee] <= 32'h34796214 ;
    mem[8'hef] <= 32'hb51eb461 ;
    mem[8'hf0] <= 32'h1625fe6f ;
    mem[8'hf1] <= 32'h9742281a ;
    mem[8'hf2] <= 32'h102b4f32 ;
    mem[8'hf3] <= 32'h914c9947 ;
    mem[8'hf4] <= 32'h1a389cd5 ;
    mem[8'hf5] <= 32'h9b5f4aa0 ;
    mem[8'hf6] <= 32'h1c362d88 ;
    mem[8'hf7] <= 32'h9d51fbfd ;
    mem[8'hf8] <= 32'he1f3b1b ;
    mem[8'hf9] <= 32'h8f78ed6e ;
    mem[8'hfa] <= 32'h8118a46 ;
    mem[8'hfb] <= 32'h89765c33 ;
    mem[8'hfc] <= 32'h20259a1 ;
    mem[8'hfd] <= 32'h83658fd4 ;
    mem[8'hfe] <= 32'h40ce8fc ;
    mem[8'hff] <= 32'h856b3e89 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
