module crctab_ev25
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'he013a34a ;
    mem[8'h2] <= 32'hc4e65b23 ;
    mem[8'h3] <= 32'h24f5f869 ;
    mem[8'h4] <= 32'h8d0dabf1 ;
    mem[8'h5] <= 32'h6d1e08bb ;
    mem[8'h6] <= 32'h49ebf0d2 ;
    mem[8'h7] <= 32'ha9f85398 ;
    mem[8'h8] <= 32'h1eda4a55 ;
    mem[8'h9] <= 32'hfec9e91f ;
    mem[8'ha] <= 32'hda3c1176 ;
    mem[8'hb] <= 32'h3a2fb23c ;
    mem[8'hc] <= 32'h93d7e1a4 ;
    mem[8'hd] <= 32'h73c442ee ;
    mem[8'he] <= 32'h5731ba87 ;
    mem[8'hf] <= 32'hb72219cd ;
    mem[8'h10] <= 32'h3db494aa ;
    mem[8'h11] <= 32'hdda737e0 ;
    mem[8'h12] <= 32'hf952cf89 ;
    mem[8'h13] <= 32'h19416cc3 ;
    mem[8'h14] <= 32'hb0b93f5b ;
    mem[8'h15] <= 32'h50aa9c11 ;
    mem[8'h16] <= 32'h745f6478 ;
    mem[8'h17] <= 32'h944cc732 ;
    mem[8'h18] <= 32'h236edeff ;
    mem[8'h19] <= 32'hc37d7db5 ;
    mem[8'h1a] <= 32'he78885dc ;
    mem[8'h1b] <= 32'h79b2696 ;
    mem[8'h1c] <= 32'hae63750e ;
    mem[8'h1d] <= 32'h4e70d644 ;
    mem[8'h1e] <= 32'h6a852e2d ;
    mem[8'h1f] <= 32'h8a968d67 ;
    mem[8'h20] <= 32'h7b692954 ;
    mem[8'h21] <= 32'h9b7a8a1e ;
    mem[8'h22] <= 32'hbf8f7277 ;
    mem[8'h23] <= 32'h5f9cd13d ;
    mem[8'h24] <= 32'hf66482a5 ;
    mem[8'h25] <= 32'h167721ef ;
    mem[8'h26] <= 32'h3282d986 ;
    mem[8'h27] <= 32'hd2917acc ;
    mem[8'h28] <= 32'h65b36301 ;
    mem[8'h29] <= 32'h85a0c04b ;
    mem[8'h2a] <= 32'ha1553822 ;
    mem[8'h2b] <= 32'h41469b68 ;
    mem[8'h2c] <= 32'he8bec8f0 ;
    mem[8'h2d] <= 32'h8ad6bba ;
    mem[8'h2e] <= 32'h2c5893d3 ;
    mem[8'h2f] <= 32'hcc4b3099 ;
    mem[8'h30] <= 32'h46ddbdfe ;
    mem[8'h31] <= 32'ha6ce1eb4 ;
    mem[8'h32] <= 32'h823be6dd ;
    mem[8'h33] <= 32'h62284597 ;
    mem[8'h34] <= 32'hcbd0160f ;
    mem[8'h35] <= 32'h2bc3b545 ;
    mem[8'h36] <= 32'hf364d2c ;
    mem[8'h37] <= 32'hef25ee66 ;
    mem[8'h38] <= 32'h5807f7ab ;
    mem[8'h39] <= 32'hb81454e1 ;
    mem[8'h3a] <= 32'h9ce1ac88 ;
    mem[8'h3b] <= 32'h7cf20fc2 ;
    mem[8'h3c] <= 32'hd50a5c5a ;
    mem[8'h3d] <= 32'h3519ff10 ;
    mem[8'h3e] <= 32'h11ec0779 ;
    mem[8'h3f] <= 32'hf1ffa433 ;
    mem[8'h40] <= 32'hf6d252a8 ;
    mem[8'h41] <= 32'h16c1f1e2 ;
    mem[8'h42] <= 32'h3234098b ;
    mem[8'h43] <= 32'hd227aac1 ;
    mem[8'h44] <= 32'h7bdff959 ;
    mem[8'h45] <= 32'h9bcc5a13 ;
    mem[8'h46] <= 32'hbf39a27a ;
    mem[8'h47] <= 32'h5f2a0130 ;
    mem[8'h48] <= 32'he80818fd ;
    mem[8'h49] <= 32'h81bbbb7 ;
    mem[8'h4a] <= 32'h2cee43de ;
    mem[8'h4b] <= 32'hccfde094 ;
    mem[8'h4c] <= 32'h6505b30c ;
    mem[8'h4d] <= 32'h85161046 ;
    mem[8'h4e] <= 32'ha1e3e82f ;
    mem[8'h4f] <= 32'h41f04b65 ;
    mem[8'h50] <= 32'hcb66c602 ;
    mem[8'h51] <= 32'h2b756548 ;
    mem[8'h52] <= 32'hf809d21 ;
    mem[8'h53] <= 32'hef933e6b ;
    mem[8'h54] <= 32'h466b6df3 ;
    mem[8'h55] <= 32'ha678ceb9 ;
    mem[8'h56] <= 32'h828d36d0 ;
    mem[8'h57] <= 32'h629e959a ;
    mem[8'h58] <= 32'hd5bc8c57 ;
    mem[8'h59] <= 32'h35af2f1d ;
    mem[8'h5a] <= 32'h115ad774 ;
    mem[8'h5b] <= 32'hf149743e ;
    mem[8'h5c] <= 32'h58b127a6 ;
    mem[8'h5d] <= 32'hb8a284ec ;
    mem[8'h5e] <= 32'h9c577c85 ;
    mem[8'h5f] <= 32'h7c44dfcf ;
    mem[8'h60] <= 32'h8dbb7bfc ;
    mem[8'h61] <= 32'h6da8d8b6 ;
    mem[8'h62] <= 32'h495d20df ;
    mem[8'h63] <= 32'ha94e8395 ;
    mem[8'h64] <= 32'hb6d00d ;
    mem[8'h65] <= 32'he0a57347 ;
    mem[8'h66] <= 32'hc4508b2e ;
    mem[8'h67] <= 32'h24432864 ;
    mem[8'h68] <= 32'h936131a9 ;
    mem[8'h69] <= 32'h737292e3 ;
    mem[8'h6a] <= 32'h57876a8a ;
    mem[8'h6b] <= 32'hb794c9c0 ;
    mem[8'h6c] <= 32'h1e6c9a58 ;
    mem[8'h6d] <= 32'hfe7f3912 ;
    mem[8'h6e] <= 32'hda8ac17b ;
    mem[8'h6f] <= 32'h3a996231 ;
    mem[8'h70] <= 32'hb00fef56 ;
    mem[8'h71] <= 32'h501c4c1c ;
    mem[8'h72] <= 32'h74e9b475 ;
    mem[8'h73] <= 32'h94fa173f ;
    mem[8'h74] <= 32'h3d0244a7 ;
    mem[8'h75] <= 32'hdd11e7ed ;
    mem[8'h76] <= 32'hf9e41f84 ;
    mem[8'h77] <= 32'h19f7bcce ;
    mem[8'h78] <= 32'haed5a503 ;
    mem[8'h79] <= 32'h4ec60649 ;
    mem[8'h7a] <= 32'h6a33fe20 ;
    mem[8'h7b] <= 32'h8a205d6a ;
    mem[8'h7c] <= 32'h23d80ef2 ;
    mem[8'h7d] <= 32'hc3cbadb8 ;
    mem[8'h7e] <= 32'he73e55d1 ;
    mem[8'h7f] <= 32'h72df69b ;
    mem[8'h80] <= 32'he965b8e7 ;
    mem[8'h81] <= 32'h9761bad ;
    mem[8'h82] <= 32'h2d83e3c4 ;
    mem[8'h83] <= 32'hcd90408e ;
    mem[8'h84] <= 32'h64681316 ;
    mem[8'h85] <= 32'h847bb05c ;
    mem[8'h86] <= 32'ha08e4835 ;
    mem[8'h87] <= 32'h409deb7f ;
    mem[8'h88] <= 32'hf7bff2b2 ;
    mem[8'h89] <= 32'h17ac51f8 ;
    mem[8'h8a] <= 32'h3359a991 ;
    mem[8'h8b] <= 32'hd34a0adb ;
    mem[8'h8c] <= 32'h7ab25943 ;
    mem[8'h8d] <= 32'h9aa1fa09 ;
    mem[8'h8e] <= 32'hbe540260 ;
    mem[8'h8f] <= 32'h5e47a12a ;
    mem[8'h90] <= 32'hd4d12c4d ;
    mem[8'h91] <= 32'h34c28f07 ;
    mem[8'h92] <= 32'h1037776e ;
    mem[8'h93] <= 32'hf024d424 ;
    mem[8'h94] <= 32'h59dc87bc ;
    mem[8'h95] <= 32'hb9cf24f6 ;
    mem[8'h96] <= 32'h9d3adc9f ;
    mem[8'h97] <= 32'h7d297fd5 ;
    mem[8'h98] <= 32'hca0b6618 ;
    mem[8'h99] <= 32'h2a18c552 ;
    mem[8'h9a] <= 32'heed3d3b ;
    mem[8'h9b] <= 32'heefe9e71 ;
    mem[8'h9c] <= 32'h4706cde9 ;
    mem[8'h9d] <= 32'ha7156ea3 ;
    mem[8'h9e] <= 32'h83e096ca ;
    mem[8'h9f] <= 32'h63f33580 ;
    mem[8'ha0] <= 32'h920c91b3 ;
    mem[8'ha1] <= 32'h721f32f9 ;
    mem[8'ha2] <= 32'h56eaca90 ;
    mem[8'ha3] <= 32'hb6f969da ;
    mem[8'ha4] <= 32'h1f013a42 ;
    mem[8'ha5] <= 32'hff129908 ;
    mem[8'ha6] <= 32'hdbe76161 ;
    mem[8'ha7] <= 32'h3bf4c22b ;
    mem[8'ha8] <= 32'h8cd6dbe6 ;
    mem[8'ha9] <= 32'h6cc578ac ;
    mem[8'haa] <= 32'h483080c5 ;
    mem[8'hab] <= 32'ha823238f ;
    mem[8'hac] <= 32'h1db7017 ;
    mem[8'had] <= 32'he1c8d35d ;
    mem[8'hae] <= 32'hc53d2b34 ;
    mem[8'haf] <= 32'h252e887e ;
    mem[8'hb0] <= 32'hafb80519 ;
    mem[8'hb1] <= 32'h4faba653 ;
    mem[8'hb2] <= 32'h6b5e5e3a ;
    mem[8'hb3] <= 32'h8b4dfd70 ;
    mem[8'hb4] <= 32'h22b5aee8 ;
    mem[8'hb5] <= 32'hc2a60da2 ;
    mem[8'hb6] <= 32'he653f5cb ;
    mem[8'hb7] <= 32'h6405681 ;
    mem[8'hb8] <= 32'hb1624f4c ;
    mem[8'hb9] <= 32'h5171ec06 ;
    mem[8'hba] <= 32'h7584146f ;
    mem[8'hbb] <= 32'h9597b725 ;
    mem[8'hbc] <= 32'h3c6fe4bd ;
    mem[8'hbd] <= 32'hdc7c47f7 ;
    mem[8'hbe] <= 32'hf889bf9e ;
    mem[8'hbf] <= 32'h189a1cd4 ;
    mem[8'hc0] <= 32'h1fb7ea4f ;
    mem[8'hc1] <= 32'hffa44905 ;
    mem[8'hc2] <= 32'hdb51b16c ;
    mem[8'hc3] <= 32'h3b421226 ;
    mem[8'hc4] <= 32'h92ba41be ;
    mem[8'hc5] <= 32'h72a9e2f4 ;
    mem[8'hc6] <= 32'h565c1a9d ;
    mem[8'hc7] <= 32'hb64fb9d7 ;
    mem[8'hc8] <= 32'h16da01a ;
    mem[8'hc9] <= 32'he17e0350 ;
    mem[8'hca] <= 32'hc58bfb39 ;
    mem[8'hcb] <= 32'h25985873 ;
    mem[8'hcc] <= 32'h8c600beb ;
    mem[8'hcd] <= 32'h6c73a8a1 ;
    mem[8'hce] <= 32'h488650c8 ;
    mem[8'hcf] <= 32'ha895f382 ;
    mem[8'hd0] <= 32'h22037ee5 ;
    mem[8'hd1] <= 32'hc210ddaf ;
    mem[8'hd2] <= 32'he6e525c6 ;
    mem[8'hd3] <= 32'h6f6868c ;
    mem[8'hd4] <= 32'haf0ed514 ;
    mem[8'hd5] <= 32'h4f1d765e ;
    mem[8'hd6] <= 32'h6be88e37 ;
    mem[8'hd7] <= 32'h8bfb2d7d ;
    mem[8'hd8] <= 32'h3cd934b0 ;
    mem[8'hd9] <= 32'hdcca97fa ;
    mem[8'hda] <= 32'hf83f6f93 ;
    mem[8'hdb] <= 32'h182cccd9 ;
    mem[8'hdc] <= 32'hb1d49f41 ;
    mem[8'hdd] <= 32'h51c73c0b ;
    mem[8'hde] <= 32'h7532c462 ;
    mem[8'hdf] <= 32'h95216728 ;
    mem[8'he0] <= 32'h64dec31b ;
    mem[8'he1] <= 32'h84cd6051 ;
    mem[8'he2] <= 32'ha0389838 ;
    mem[8'he3] <= 32'h402b3b72 ;
    mem[8'he4] <= 32'he9d368ea ;
    mem[8'he5] <= 32'h9c0cba0 ;
    mem[8'he6] <= 32'h2d3533c9 ;
    mem[8'he7] <= 32'hcd269083 ;
    mem[8'he8] <= 32'h7a04894e ;
    mem[8'he9] <= 32'h9a172a04 ;
    mem[8'hea] <= 32'hbee2d26d ;
    mem[8'heb] <= 32'h5ef17127 ;
    mem[8'hec] <= 32'hf70922bf ;
    mem[8'hed] <= 32'h171a81f5 ;
    mem[8'hee] <= 32'h33ef799c ;
    mem[8'hef] <= 32'hd3fcdad6 ;
    mem[8'hf0] <= 32'h596a57b1 ;
    mem[8'hf1] <= 32'hb979f4fb ;
    mem[8'hf2] <= 32'h9d8c0c92 ;
    mem[8'hf3] <= 32'h7d9fafd8 ;
    mem[8'hf4] <= 32'hd467fc40 ;
    mem[8'hf5] <= 32'h34745f0a ;
    mem[8'hf6] <= 32'h1081a763 ;
    mem[8'hf7] <= 32'hf0920429 ;
    mem[8'hf8] <= 32'h47b01de4 ;
    mem[8'hf9] <= 32'ha7a3beae ;
    mem[8'hfa] <= 32'h835646c7 ;
    mem[8'hfb] <= 32'h6345e58d ;
    mem[8'hfc] <= 32'hcabdb615 ;
    mem[8'hfd] <= 32'h2aae155f ;
    mem[8'hfe] <= 32'he5bed36 ;
    mem[8'hff] <= 32'hee484e7c ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
