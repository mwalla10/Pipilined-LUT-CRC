module crctab_ev16
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h17d3315d ;
    mem[8'h2] <= 32'h2fa662ba ;
    mem[8'h3] <= 32'h387553e7 ;
    mem[8'h4] <= 32'h5f4cc574 ;
    mem[8'h5] <= 32'h489ff429 ;
    mem[8'h6] <= 32'h70eaa7ce ;
    mem[8'h7] <= 32'h67399693 ;
    mem[8'h8] <= 32'hbe998ae8 ;
    mem[8'h9] <= 32'ha94abbb5 ;
    mem[8'ha] <= 32'h913fe852 ;
    mem[8'hb] <= 32'h86ecd90f ;
    mem[8'hc] <= 32'he1d54f9c ;
    mem[8'hd] <= 32'hf6067ec1 ;
    mem[8'he] <= 32'hce732d26 ;
    mem[8'hf] <= 32'hd9a01c7b ;
    mem[8'h10] <= 32'h79f20867 ;
    mem[8'h11] <= 32'h6e21393a ;
    mem[8'h12] <= 32'h56546add ;
    mem[8'h13] <= 32'h41875b80 ;
    mem[8'h14] <= 32'h26becd13 ;
    mem[8'h15] <= 32'h316dfc4e ;
    mem[8'h16] <= 32'h918afa9 ;
    mem[8'h17] <= 32'h1ecb9ef4 ;
    mem[8'h18] <= 32'hc76b828f ;
    mem[8'h19] <= 32'hd0b8b3d2 ;
    mem[8'h1a] <= 32'he8cde035 ;
    mem[8'h1b] <= 32'hff1ed168 ;
    mem[8'h1c] <= 32'h982747fb ;
    mem[8'h1d] <= 32'h8ff476a6 ;
    mem[8'h1e] <= 32'hb7812541 ;
    mem[8'h1f] <= 32'ha052141c ;
    mem[8'h20] <= 32'hf3e410ce ;
    mem[8'h21] <= 32'he4372193 ;
    mem[8'h22] <= 32'hdc427274 ;
    mem[8'h23] <= 32'hcb914329 ;
    mem[8'h24] <= 32'haca8d5ba ;
    mem[8'h25] <= 32'hbb7be4e7 ;
    mem[8'h26] <= 32'h830eb700 ;
    mem[8'h27] <= 32'h94dd865d ;
    mem[8'h28] <= 32'h4d7d9a26 ;
    mem[8'h29] <= 32'h5aaeab7b ;
    mem[8'h2a] <= 32'h62dbf89c ;
    mem[8'h2b] <= 32'h7508c9c1 ;
    mem[8'h2c] <= 32'h12315f52 ;
    mem[8'h2d] <= 32'h5e26e0f ;
    mem[8'h2e] <= 32'h3d973de8 ;
    mem[8'h2f] <= 32'h2a440cb5 ;
    mem[8'h30] <= 32'h8a1618a9 ;
    mem[8'h31] <= 32'h9dc529f4 ;
    mem[8'h32] <= 32'ha5b07a13 ;
    mem[8'h33] <= 32'hb2634b4e ;
    mem[8'h34] <= 32'hd55adddd ;
    mem[8'h35] <= 32'hc289ec80 ;
    mem[8'h36] <= 32'hfafcbf67 ;
    mem[8'h37] <= 32'hed2f8e3a ;
    mem[8'h38] <= 32'h348f9241 ;
    mem[8'h39] <= 32'h235ca31c ;
    mem[8'h3a] <= 32'h1b29f0fb ;
    mem[8'h3b] <= 32'hcfac1a6 ;
    mem[8'h3c] <= 32'h6bc35735 ;
    mem[8'h3d] <= 32'h7c106668 ;
    mem[8'h3e] <= 32'h4465358f ;
    mem[8'h3f] <= 32'h53b604d2 ;
    mem[8'h40] <= 32'he3093c2b ;
    mem[8'h41] <= 32'hf4da0d76 ;
    mem[8'h42] <= 32'hccaf5e91 ;
    mem[8'h43] <= 32'hdb7c6fcc ;
    mem[8'h44] <= 32'hbc45f95f ;
    mem[8'h45] <= 32'hab96c802 ;
    mem[8'h46] <= 32'h93e39be5 ;
    mem[8'h47] <= 32'h8430aab8 ;
    mem[8'h48] <= 32'h5d90b6c3 ;
    mem[8'h49] <= 32'h4a43879e ;
    mem[8'h4a] <= 32'h7236d479 ;
    mem[8'h4b] <= 32'h65e5e524 ;
    mem[8'h4c] <= 32'h2dc73b7 ;
    mem[8'h4d] <= 32'h150f42ea ;
    mem[8'h4e] <= 32'h2d7a110d ;
    mem[8'h4f] <= 32'h3aa92050 ;
    mem[8'h50] <= 32'h9afb344c ;
    mem[8'h51] <= 32'h8d280511 ;
    mem[8'h52] <= 32'hb55d56f6 ;
    mem[8'h53] <= 32'ha28e67ab ;
    mem[8'h54] <= 32'hc5b7f138 ;
    mem[8'h55] <= 32'hd264c065 ;
    mem[8'h56] <= 32'hea119382 ;
    mem[8'h57] <= 32'hfdc2a2df ;
    mem[8'h58] <= 32'h2462bea4 ;
    mem[8'h59] <= 32'h33b18ff9 ;
    mem[8'h5a] <= 32'hbc4dc1e ;
    mem[8'h5b] <= 32'h1c17ed43 ;
    mem[8'h5c] <= 32'h7b2e7bd0 ;
    mem[8'h5d] <= 32'h6cfd4a8d ;
    mem[8'h5e] <= 32'h5488196a ;
    mem[8'h5f] <= 32'h435b2837 ;
    mem[8'h60] <= 32'h10ed2ce5 ;
    mem[8'h61] <= 32'h73e1db8 ;
    mem[8'h62] <= 32'h3f4b4e5f ;
    mem[8'h63] <= 32'h28987f02 ;
    mem[8'h64] <= 32'h4fa1e991 ;
    mem[8'h65] <= 32'h5872d8cc ;
    mem[8'h66] <= 32'h60078b2b ;
    mem[8'h67] <= 32'h77d4ba76 ;
    mem[8'h68] <= 32'hae74a60d ;
    mem[8'h69] <= 32'hb9a79750 ;
    mem[8'h6a] <= 32'h81d2c4b7 ;
    mem[8'h6b] <= 32'h9601f5ea ;
    mem[8'h6c] <= 32'hf1386379 ;
    mem[8'h6d] <= 32'he6eb5224 ;
    mem[8'h6e] <= 32'hde9e01c3 ;
    mem[8'h6f] <= 32'hc94d309e ;
    mem[8'h70] <= 32'h691f2482 ;
    mem[8'h71] <= 32'h7ecc15df ;
    mem[8'h72] <= 32'h46b94638 ;
    mem[8'h73] <= 32'h516a7765 ;
    mem[8'h74] <= 32'h3653e1f6 ;
    mem[8'h75] <= 32'h2180d0ab ;
    mem[8'h76] <= 32'h19f5834c ;
    mem[8'h77] <= 32'he26b211 ;
    mem[8'h78] <= 32'hd786ae6a ;
    mem[8'h79] <= 32'hc0559f37 ;
    mem[8'h7a] <= 32'hf820ccd0 ;
    mem[8'h7b] <= 32'heff3fd8d ;
    mem[8'h7c] <= 32'h88ca6b1e ;
    mem[8'h7d] <= 32'h9f195a43 ;
    mem[8'h7e] <= 32'ha76c09a4 ;
    mem[8'h7f] <= 32'hb0bf38f9 ;
    mem[8'h80] <= 32'hc2d365e1 ;
    mem[8'h81] <= 32'hd50054bc ;
    mem[8'h82] <= 32'hed75075b ;
    mem[8'h83] <= 32'hfaa63606 ;
    mem[8'h84] <= 32'h9d9fa095 ;
    mem[8'h85] <= 32'h8a4c91c8 ;
    mem[8'h86] <= 32'hb239c22f ;
    mem[8'h87] <= 32'ha5eaf372 ;
    mem[8'h88] <= 32'h7c4aef09 ;
    mem[8'h89] <= 32'h6b99de54 ;
    mem[8'h8a] <= 32'h53ec8db3 ;
    mem[8'h8b] <= 32'h443fbcee ;
    mem[8'h8c] <= 32'h23062a7d ;
    mem[8'h8d] <= 32'h34d51b20 ;
    mem[8'h8e] <= 32'hca048c7 ;
    mem[8'h8f] <= 32'h1b73799a ;
    mem[8'h90] <= 32'hbb216d86 ;
    mem[8'h91] <= 32'hacf25cdb ;
    mem[8'h92] <= 32'h94870f3c ;
    mem[8'h93] <= 32'h83543e61 ;
    mem[8'h94] <= 32'he46da8f2 ;
    mem[8'h95] <= 32'hf3be99af ;
    mem[8'h96] <= 32'hcbcbca48 ;
    mem[8'h97] <= 32'hdc18fb15 ;
    mem[8'h98] <= 32'h5b8e76e ;
    mem[8'h99] <= 32'h126bd633 ;
    mem[8'h9a] <= 32'h2a1e85d4 ;
    mem[8'h9b] <= 32'h3dcdb489 ;
    mem[8'h9c] <= 32'h5af4221a ;
    mem[8'h9d] <= 32'h4d271347 ;
    mem[8'h9e] <= 32'h755240a0 ;
    mem[8'h9f] <= 32'h628171fd ;
    mem[8'ha0] <= 32'h3137752f ;
    mem[8'ha1] <= 32'h26e44472 ;
    mem[8'ha2] <= 32'h1e911795 ;
    mem[8'ha3] <= 32'h94226c8 ;
    mem[8'ha4] <= 32'h6e7bb05b ;
    mem[8'ha5] <= 32'h79a88106 ;
    mem[8'ha6] <= 32'h41ddd2e1 ;
    mem[8'ha7] <= 32'h560ee3bc ;
    mem[8'ha8] <= 32'h8faeffc7 ;
    mem[8'ha9] <= 32'h987dce9a ;
    mem[8'haa] <= 32'ha0089d7d ;
    mem[8'hab] <= 32'hb7dbac20 ;
    mem[8'hac] <= 32'hd0e23ab3 ;
    mem[8'had] <= 32'hc7310bee ;
    mem[8'hae] <= 32'hff445809 ;
    mem[8'haf] <= 32'he8976954 ;
    mem[8'hb0] <= 32'h48c57d48 ;
    mem[8'hb1] <= 32'h5f164c15 ;
    mem[8'hb2] <= 32'h67631ff2 ;
    mem[8'hb3] <= 32'h70b02eaf ;
    mem[8'hb4] <= 32'h1789b83c ;
    mem[8'hb5] <= 32'h5a8961 ;
    mem[8'hb6] <= 32'h382fda86 ;
    mem[8'hb7] <= 32'h2ffcebdb ;
    mem[8'hb8] <= 32'hf65cf7a0 ;
    mem[8'hb9] <= 32'he18fc6fd ;
    mem[8'hba] <= 32'hd9fa951a ;
    mem[8'hbb] <= 32'hce29a447 ;
    mem[8'hbc] <= 32'ha91032d4 ;
    mem[8'hbd] <= 32'hbec30389 ;
    mem[8'hbe] <= 32'h86b6506e ;
    mem[8'hbf] <= 32'h91656133 ;
    mem[8'hc0] <= 32'h21da59ca ;
    mem[8'hc1] <= 32'h36096897 ;
    mem[8'hc2] <= 32'he7c3b70 ;
    mem[8'hc3] <= 32'h19af0a2d ;
    mem[8'hc4] <= 32'h7e969cbe ;
    mem[8'hc5] <= 32'h6945ade3 ;
    mem[8'hc6] <= 32'h5130fe04 ;
    mem[8'hc7] <= 32'h46e3cf59 ;
    mem[8'hc8] <= 32'h9f43d322 ;
    mem[8'hc9] <= 32'h8890e27f ;
    mem[8'hca] <= 32'hb0e5b198 ;
    mem[8'hcb] <= 32'ha73680c5 ;
    mem[8'hcc] <= 32'hc00f1656 ;
    mem[8'hcd] <= 32'hd7dc270b ;
    mem[8'hce] <= 32'hefa974ec ;
    mem[8'hcf] <= 32'hf87a45b1 ;
    mem[8'hd0] <= 32'h582851ad ;
    mem[8'hd1] <= 32'h4ffb60f0 ;
    mem[8'hd2] <= 32'h778e3317 ;
    mem[8'hd3] <= 32'h605d024a ;
    mem[8'hd4] <= 32'h76494d9 ;
    mem[8'hd5] <= 32'h10b7a584 ;
    mem[8'hd6] <= 32'h28c2f663 ;
    mem[8'hd7] <= 32'h3f11c73e ;
    mem[8'hd8] <= 32'he6b1db45 ;
    mem[8'hd9] <= 32'hf162ea18 ;
    mem[8'hda] <= 32'hc917b9ff ;
    mem[8'hdb] <= 32'hdec488a2 ;
    mem[8'hdc] <= 32'hb9fd1e31 ;
    mem[8'hdd] <= 32'hae2e2f6c ;
    mem[8'hde] <= 32'h965b7c8b ;
    mem[8'hdf] <= 32'h81884dd6 ;
    mem[8'he0] <= 32'hd23e4904 ;
    mem[8'he1] <= 32'hc5ed7859 ;
    mem[8'he2] <= 32'hfd982bbe ;
    mem[8'he3] <= 32'hea4b1ae3 ;
    mem[8'he4] <= 32'h8d728c70 ;
    mem[8'he5] <= 32'h9aa1bd2d ;
    mem[8'he6] <= 32'ha2d4eeca ;
    mem[8'he7] <= 32'hb507df97 ;
    mem[8'he8] <= 32'h6ca7c3ec ;
    mem[8'he9] <= 32'h7b74f2b1 ;
    mem[8'hea] <= 32'h4301a156 ;
    mem[8'heb] <= 32'h54d2900b ;
    mem[8'hec] <= 32'h33eb0698 ;
    mem[8'hed] <= 32'h243837c5 ;
    mem[8'hee] <= 32'h1c4d6422 ;
    mem[8'hef] <= 32'hb9e557f ;
    mem[8'hf0] <= 32'habcc4163 ;
    mem[8'hf1] <= 32'hbc1f703e ;
    mem[8'hf2] <= 32'h846a23d9 ;
    mem[8'hf3] <= 32'h93b91284 ;
    mem[8'hf4] <= 32'hf4808417 ;
    mem[8'hf5] <= 32'he353b54a ;
    mem[8'hf6] <= 32'hdb26e6ad ;
    mem[8'hf7] <= 32'hccf5d7f0 ;
    mem[8'hf8] <= 32'h1555cb8b ;
    mem[8'hf9] <= 32'h286fad6 ;
    mem[8'hfa] <= 32'h3af3a931 ;
    mem[8'hfb] <= 32'h2d20986c ;
    mem[8'hfc] <= 32'h4a190eff ;
    mem[8'hfd] <= 32'h5dca3fa2 ;
    mem[8'hfe] <= 32'h65bf6c45 ;
    mem[8'hff] <= 32'h726c5d18 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
