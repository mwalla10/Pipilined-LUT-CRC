module crctab_ev20
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'hc5b9cd4c ;
    mem[8'h2] <= 32'h8fb2872f ;
    mem[8'h3] <= 32'h4a0b4a63 ;
    mem[8'h4] <= 32'h1ba413e9 ;
    mem[8'h5] <= 32'hde1ddea5 ;
    mem[8'h6] <= 32'h941694c6 ;
    mem[8'h7] <= 32'h51af598a ;
    mem[8'h8] <= 32'h374827d2 ;
    mem[8'h9] <= 32'hf2f1ea9e ;
    mem[8'ha] <= 32'hb8faa0fd ;
    mem[8'hb] <= 32'h7d436db1 ;
    mem[8'hc] <= 32'h2cec343b ;
    mem[8'hd] <= 32'he955f977 ;
    mem[8'he] <= 32'ha35eb314 ;
    mem[8'hf] <= 32'h66e77e58 ;
    mem[8'h10] <= 32'h6e904fa4 ;
    mem[8'h11] <= 32'hab2982e8 ;
    mem[8'h12] <= 32'he122c88b ;
    mem[8'h13] <= 32'h249b05c7 ;
    mem[8'h14] <= 32'h75345c4d ;
    mem[8'h15] <= 32'hb08d9101 ;
    mem[8'h16] <= 32'hfa86db62 ;
    mem[8'h17] <= 32'h3f3f162e ;
    mem[8'h18] <= 32'h59d86876 ;
    mem[8'h19] <= 32'h9c61a53a ;
    mem[8'h1a] <= 32'hd66aef59 ;
    mem[8'h1b] <= 32'h13d32215 ;
    mem[8'h1c] <= 32'h427c7b9f ;
    mem[8'h1d] <= 32'h87c5b6d3 ;
    mem[8'h1e] <= 32'hcdcefcb0 ;
    mem[8'h1f] <= 32'h87731fc ;
    mem[8'h20] <= 32'hdd209f48 ;
    mem[8'h21] <= 32'h18995204 ;
    mem[8'h22] <= 32'h52921867 ;
    mem[8'h23] <= 32'h972bd52b ;
    mem[8'h24] <= 32'hc6848ca1 ;
    mem[8'h25] <= 32'h33d41ed ;
    mem[8'h26] <= 32'h49360b8e ;
    mem[8'h27] <= 32'h8c8fc6c2 ;
    mem[8'h28] <= 32'hea68b89a ;
    mem[8'h29] <= 32'h2fd175d6 ;
    mem[8'h2a] <= 32'h65da3fb5 ;
    mem[8'h2b] <= 32'ha063f2f9 ;
    mem[8'h2c] <= 32'hf1ccab73 ;
    mem[8'h2d] <= 32'h3475663f ;
    mem[8'h2e] <= 32'h7e7e2c5c ;
    mem[8'h2f] <= 32'hbbc7e110 ;
    mem[8'h30] <= 32'hb3b0d0ec ;
    mem[8'h31] <= 32'h76091da0 ;
    mem[8'h32] <= 32'h3c0257c3 ;
    mem[8'h33] <= 32'hf9bb9a8f ;
    mem[8'h34] <= 32'ha814c305 ;
    mem[8'h35] <= 32'h6dad0e49 ;
    mem[8'h36] <= 32'h27a6442a ;
    mem[8'h37] <= 32'he21f8966 ;
    mem[8'h38] <= 32'h84f8f73e ;
    mem[8'h39] <= 32'h41413a72 ;
    mem[8'h3a] <= 32'hb4a7011 ;
    mem[8'h3b] <= 32'hcef3bd5d ;
    mem[8'h3c] <= 32'h9f5ce4d7 ;
    mem[8'h3d] <= 32'h5ae5299b ;
    mem[8'h3e] <= 32'h10ee63f8 ;
    mem[8'h3f] <= 32'hd557aeb4 ;
    mem[8'h40] <= 32'hbe802327 ;
    mem[8'h41] <= 32'h7b39ee6b ;
    mem[8'h42] <= 32'h3132a408 ;
    mem[8'h43] <= 32'hf48b6944 ;
    mem[8'h44] <= 32'ha52430ce ;
    mem[8'h45] <= 32'h609dfd82 ;
    mem[8'h46] <= 32'h2a96b7e1 ;
    mem[8'h47] <= 32'hef2f7aad ;
    mem[8'h48] <= 32'h89c804f5 ;
    mem[8'h49] <= 32'h4c71c9b9 ;
    mem[8'h4a] <= 32'h67a83da ;
    mem[8'h4b] <= 32'hc3c34e96 ;
    mem[8'h4c] <= 32'h926c171c ;
    mem[8'h4d] <= 32'h57d5da50 ;
    mem[8'h4e] <= 32'h1dde9033 ;
    mem[8'h4f] <= 32'hd8675d7f ;
    mem[8'h50] <= 32'hd0106c83 ;
    mem[8'h51] <= 32'h15a9a1cf ;
    mem[8'h52] <= 32'h5fa2ebac ;
    mem[8'h53] <= 32'h9a1b26e0 ;
    mem[8'h54] <= 32'hcbb47f6a ;
    mem[8'h55] <= 32'he0db226 ;
    mem[8'h56] <= 32'h4406f845 ;
    mem[8'h57] <= 32'h81bf3509 ;
    mem[8'h58] <= 32'he7584b51 ;
    mem[8'h59] <= 32'h22e1861d ;
    mem[8'h5a] <= 32'h68eacc7e ;
    mem[8'h5b] <= 32'had530132 ;
    mem[8'h5c] <= 32'hfcfc58b8 ;
    mem[8'h5d] <= 32'h394595f4 ;
    mem[8'h5e] <= 32'h734edf97 ;
    mem[8'h5f] <= 32'hb6f712db ;
    mem[8'h60] <= 32'h63a0bc6f ;
    mem[8'h61] <= 32'ha6197123 ;
    mem[8'h62] <= 32'hec123b40 ;
    mem[8'h63] <= 32'h29abf60c ;
    mem[8'h64] <= 32'h7804af86 ;
    mem[8'h65] <= 32'hbdbd62ca ;
    mem[8'h66] <= 32'hf7b628a9 ;
    mem[8'h67] <= 32'h320fe5e5 ;
    mem[8'h68] <= 32'h54e89bbd ;
    mem[8'h69] <= 32'h915156f1 ;
    mem[8'h6a] <= 32'hdb5a1c92 ;
    mem[8'h6b] <= 32'h1ee3d1de ;
    mem[8'h6c] <= 32'h4f4c8854 ;
    mem[8'h6d] <= 32'h8af54518 ;
    mem[8'h6e] <= 32'hc0fe0f7b ;
    mem[8'h6f] <= 32'h547c237 ;
    mem[8'h70] <= 32'hd30f3cb ;
    mem[8'h71] <= 32'hc8893e87 ;
    mem[8'h72] <= 32'h828274e4 ;
    mem[8'h73] <= 32'h473bb9a8 ;
    mem[8'h74] <= 32'h1694e022 ;
    mem[8'h75] <= 32'hd32d2d6e ;
    mem[8'h76] <= 32'h9926670d ;
    mem[8'h77] <= 32'h5c9faa41 ;
    mem[8'h78] <= 32'h3a78d419 ;
    mem[8'h79] <= 32'hffc11955 ;
    mem[8'h7a] <= 32'hb5ca5336 ;
    mem[8'h7b] <= 32'h70739e7a ;
    mem[8'h7c] <= 32'h21dcc7f0 ;
    mem[8'h7d] <= 32'he4650abc ;
    mem[8'h7e] <= 32'hae6e40df ;
    mem[8'h7f] <= 32'h6bd78d93 ;
    mem[8'h80] <= 32'h79c15bf9 ;
    mem[8'h81] <= 32'hbc7896b5 ;
    mem[8'h82] <= 32'hf673dcd6 ;
    mem[8'h83] <= 32'h33ca119a ;
    mem[8'h84] <= 32'h62654810 ;
    mem[8'h85] <= 32'ha7dc855c ;
    mem[8'h86] <= 32'hedd7cf3f ;
    mem[8'h87] <= 32'h286e0273 ;
    mem[8'h88] <= 32'h4e897c2b ;
    mem[8'h89] <= 32'h8b30b167 ;
    mem[8'h8a] <= 32'hc13bfb04 ;
    mem[8'h8b] <= 32'h4823648 ;
    mem[8'h8c] <= 32'h552d6fc2 ;
    mem[8'h8d] <= 32'h9094a28e ;
    mem[8'h8e] <= 32'hda9fe8ed ;
    mem[8'h8f] <= 32'h1f2625a1 ;
    mem[8'h90] <= 32'h1751145d ;
    mem[8'h91] <= 32'hd2e8d911 ;
    mem[8'h92] <= 32'h98e39372 ;
    mem[8'h93] <= 32'h5d5a5e3e ;
    mem[8'h94] <= 32'hcf507b4 ;
    mem[8'h95] <= 32'hc94ccaf8 ;
    mem[8'h96] <= 32'h8347809b ;
    mem[8'h97] <= 32'h46fe4dd7 ;
    mem[8'h98] <= 32'h2019338f ;
    mem[8'h99] <= 32'he5a0fec3 ;
    mem[8'h9a] <= 32'hafabb4a0 ;
    mem[8'h9b] <= 32'h6a1279ec ;
    mem[8'h9c] <= 32'h3bbd2066 ;
    mem[8'h9d] <= 32'hfe04ed2a ;
    mem[8'h9e] <= 32'hb40fa749 ;
    mem[8'h9f] <= 32'h71b66a05 ;
    mem[8'ha0] <= 32'ha4e1c4b1 ;
    mem[8'ha1] <= 32'h615809fd ;
    mem[8'ha2] <= 32'h2b53439e ;
    mem[8'ha3] <= 32'heeea8ed2 ;
    mem[8'ha4] <= 32'hbf45d758 ;
    mem[8'ha5] <= 32'h7afc1a14 ;
    mem[8'ha6] <= 32'h30f75077 ;
    mem[8'ha7] <= 32'hf54e9d3b ;
    mem[8'ha8] <= 32'h93a9e363 ;
    mem[8'ha9] <= 32'h56102e2f ;
    mem[8'haa] <= 32'h1c1b644c ;
    mem[8'hab] <= 32'hd9a2a900 ;
    mem[8'hac] <= 32'h880df08a ;
    mem[8'had] <= 32'h4db43dc6 ;
    mem[8'hae] <= 32'h7bf77a5 ;
    mem[8'haf] <= 32'hc206bae9 ;
    mem[8'hb0] <= 32'hca718b15 ;
    mem[8'hb1] <= 32'hfc84659 ;
    mem[8'hb2] <= 32'h45c30c3a ;
    mem[8'hb3] <= 32'h807ac176 ;
    mem[8'hb4] <= 32'hd1d598fc ;
    mem[8'hb5] <= 32'h146c55b0 ;
    mem[8'hb6] <= 32'h5e671fd3 ;
    mem[8'hb7] <= 32'h9bded29f ;
    mem[8'hb8] <= 32'hfd39acc7 ;
    mem[8'hb9] <= 32'h3880618b ;
    mem[8'hba] <= 32'h728b2be8 ;
    mem[8'hbb] <= 32'hb732e6a4 ;
    mem[8'hbc] <= 32'he69dbf2e ;
    mem[8'hbd] <= 32'h23247262 ;
    mem[8'hbe] <= 32'h692f3801 ;
    mem[8'hbf] <= 32'hac96f54d ;
    mem[8'hc0] <= 32'hc74178de ;
    mem[8'hc1] <= 32'h2f8b592 ;
    mem[8'hc2] <= 32'h48f3fff1 ;
    mem[8'hc3] <= 32'h8d4a32bd ;
    mem[8'hc4] <= 32'hdce56b37 ;
    mem[8'hc5] <= 32'h195ca67b ;
    mem[8'hc6] <= 32'h5357ec18 ;
    mem[8'hc7] <= 32'h96ee2154 ;
    mem[8'hc8] <= 32'hf0095f0c ;
    mem[8'hc9] <= 32'h35b09240 ;
    mem[8'hca] <= 32'h7fbbd823 ;
    mem[8'hcb] <= 32'hba02156f ;
    mem[8'hcc] <= 32'hebad4ce5 ;
    mem[8'hcd] <= 32'h2e1481a9 ;
    mem[8'hce] <= 32'h641fcbca ;
    mem[8'hcf] <= 32'ha1a60686 ;
    mem[8'hd0] <= 32'ha9d1377a ;
    mem[8'hd1] <= 32'h6c68fa36 ;
    mem[8'hd2] <= 32'h2663b055 ;
    mem[8'hd3] <= 32'he3da7d19 ;
    mem[8'hd4] <= 32'hb2752493 ;
    mem[8'hd5] <= 32'h77cce9df ;
    mem[8'hd6] <= 32'h3dc7a3bc ;
    mem[8'hd7] <= 32'hf87e6ef0 ;
    mem[8'hd8] <= 32'h9e9910a8 ;
    mem[8'hd9] <= 32'h5b20dde4 ;
    mem[8'hda] <= 32'h112b9787 ;
    mem[8'hdb] <= 32'hd4925acb ;
    mem[8'hdc] <= 32'h853d0341 ;
    mem[8'hdd] <= 32'h4084ce0d ;
    mem[8'hde] <= 32'ha8f846e ;
    mem[8'hdf] <= 32'hcf364922 ;
    mem[8'he0] <= 32'h1a61e796 ;
    mem[8'he1] <= 32'hdfd82ada ;
    mem[8'he2] <= 32'h95d360b9 ;
    mem[8'he3] <= 32'h506aadf5 ;
    mem[8'he4] <= 32'h1c5f47f ;
    mem[8'he5] <= 32'hc47c3933 ;
    mem[8'he6] <= 32'h8e777350 ;
    mem[8'he7] <= 32'h4bcebe1c ;
    mem[8'he8] <= 32'h2d29c044 ;
    mem[8'he9] <= 32'he8900d08 ;
    mem[8'hea] <= 32'ha29b476b ;
    mem[8'heb] <= 32'h67228a27 ;
    mem[8'hec] <= 32'h368dd3ad ;
    mem[8'hed] <= 32'hf3341ee1 ;
    mem[8'hee] <= 32'hb93f5482 ;
    mem[8'hef] <= 32'h7c8699ce ;
    mem[8'hf0] <= 32'h74f1a832 ;
    mem[8'hf1] <= 32'hb148657e ;
    mem[8'hf2] <= 32'hfb432f1d ;
    mem[8'hf3] <= 32'h3efae251 ;
    mem[8'hf4] <= 32'h6f55bbdb ;
    mem[8'hf5] <= 32'haaec7697 ;
    mem[8'hf6] <= 32'he0e73cf4 ;
    mem[8'hf7] <= 32'h255ef1b8 ;
    mem[8'hf8] <= 32'h43b98fe0 ;
    mem[8'hf9] <= 32'h860042ac ;
    mem[8'hfa] <= 32'hcc0b08cf ;
    mem[8'hfb] <= 32'h9b2c583 ;
    mem[8'hfc] <= 32'h581d9c09 ;
    mem[8'hfd] <= 32'h9da45145 ;
    mem[8'hfe] <= 32'hd7af1b26 ;
    mem[8'hff] <= 32'h1216d66a ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
