module crctab_ev13
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h47f7cec1 ;
    mem[8'h2] <= 32'h8fef9d82 ;
    mem[8'h3] <= 32'hc8185343 ;
    mem[8'h4] <= 32'h1b1e26b3 ;
    mem[8'h5] <= 32'h5ce9e872 ;
    mem[8'h6] <= 32'h94f1bb31 ;
    mem[8'h7] <= 32'hd30675f0 ;
    mem[8'h8] <= 32'h363c4d66 ;
    mem[8'h9] <= 32'h71cb83a7 ;
    mem[8'ha] <= 32'hb9d3d0e4 ;
    mem[8'hb] <= 32'hfe241e25 ;
    mem[8'hc] <= 32'h2d226bd5 ;
    mem[8'hd] <= 32'h6ad5a514 ;
    mem[8'he] <= 32'ha2cdf657 ;
    mem[8'hf] <= 32'he53a3896 ;
    mem[8'h10] <= 32'h6c789acc ;
    mem[8'h11] <= 32'h2b8f540d ;
    mem[8'h12] <= 32'he397074e ;
    mem[8'h13] <= 32'ha460c98f ;
    mem[8'h14] <= 32'h7766bc7f ;
    mem[8'h15] <= 32'h309172be ;
    mem[8'h16] <= 32'hf88921fd ;
    mem[8'h17] <= 32'hbf7eef3c ;
    mem[8'h18] <= 32'h5a44d7aa ;
    mem[8'h19] <= 32'h1db3196b ;
    mem[8'h1a] <= 32'hd5ab4a28 ;
    mem[8'h1b] <= 32'h925c84e9 ;
    mem[8'h1c] <= 32'h415af119 ;
    mem[8'h1d] <= 32'h6ad3fd8 ;
    mem[8'h1e] <= 32'hceb56c9b ;
    mem[8'h1f] <= 32'h8942a25a ;
    mem[8'h20] <= 32'hd8f13598 ;
    mem[8'h21] <= 32'h9f06fb59 ;
    mem[8'h22] <= 32'h571ea81a ;
    mem[8'h23] <= 32'h10e966db ;
    mem[8'h24] <= 32'hc3ef132b ;
    mem[8'h25] <= 32'h8418ddea ;
    mem[8'h26] <= 32'h4c008ea9 ;
    mem[8'h27] <= 32'hbf74068 ;
    mem[8'h28] <= 32'heecd78fe ;
    mem[8'h29] <= 32'ha93ab63f ;
    mem[8'h2a] <= 32'h6122e57c ;
    mem[8'h2b] <= 32'h26d52bbd ;
    mem[8'h2c] <= 32'hf5d35e4d ;
    mem[8'h2d] <= 32'hb224908c ;
    mem[8'h2e] <= 32'h7a3cc3cf ;
    mem[8'h2f] <= 32'h3dcb0d0e ;
    mem[8'h30] <= 32'hb489af54 ;
    mem[8'h31] <= 32'hf37e6195 ;
    mem[8'h32] <= 32'h3b6632d6 ;
    mem[8'h33] <= 32'h7c91fc17 ;
    mem[8'h34] <= 32'haf9789e7 ;
    mem[8'h35] <= 32'he8604726 ;
    mem[8'h36] <= 32'h20781465 ;
    mem[8'h37] <= 32'h678fdaa4 ;
    mem[8'h38] <= 32'h82b5e232 ;
    mem[8'h39] <= 32'hc5422cf3 ;
    mem[8'h3a] <= 32'hd5a7fb0 ;
    mem[8'h3b] <= 32'h4aadb171 ;
    mem[8'h3c] <= 32'h99abc481 ;
    mem[8'h3d] <= 32'hde5c0a40 ;
    mem[8'h3e] <= 32'h16445903 ;
    mem[8'h3f] <= 32'h51b397c2 ;
    mem[8'h40] <= 32'hb5237687 ;
    mem[8'h41] <= 32'hf2d4b846 ;
    mem[8'h42] <= 32'h3acceb05 ;
    mem[8'h43] <= 32'h7d3b25c4 ;
    mem[8'h44] <= 32'hae3d5034 ;
    mem[8'h45] <= 32'he9ca9ef5 ;
    mem[8'h46] <= 32'h21d2cdb6 ;
    mem[8'h47] <= 32'h66250377 ;
    mem[8'h48] <= 32'h831f3be1 ;
    mem[8'h49] <= 32'hc4e8f520 ;
    mem[8'h4a] <= 32'hcf0a663 ;
    mem[8'h4b] <= 32'h4b0768a2 ;
    mem[8'h4c] <= 32'h98011d52 ;
    mem[8'h4d] <= 32'hdff6d393 ;
    mem[8'h4e] <= 32'h17ee80d0 ;
    mem[8'h4f] <= 32'h50194e11 ;
    mem[8'h50] <= 32'hd95bec4b ;
    mem[8'h51] <= 32'h9eac228a ;
    mem[8'h52] <= 32'h56b471c9 ;
    mem[8'h53] <= 32'h1143bf08 ;
    mem[8'h54] <= 32'hc245caf8 ;
    mem[8'h55] <= 32'h85b20439 ;
    mem[8'h56] <= 32'h4daa577a ;
    mem[8'h57] <= 32'ha5d99bb ;
    mem[8'h58] <= 32'hef67a12d ;
    mem[8'h59] <= 32'ha8906fec ;
    mem[8'h5a] <= 32'h60883caf ;
    mem[8'h5b] <= 32'h277ff26e ;
    mem[8'h5c] <= 32'hf479879e ;
    mem[8'h5d] <= 32'hb38e495f ;
    mem[8'h5e] <= 32'h7b961a1c ;
    mem[8'h5f] <= 32'h3c61d4dd ;
    mem[8'h60] <= 32'h6dd2431f ;
    mem[8'h61] <= 32'h2a258dde ;
    mem[8'h62] <= 32'he23dde9d ;
    mem[8'h63] <= 32'ha5ca105c ;
    mem[8'h64] <= 32'h76cc65ac ;
    mem[8'h65] <= 32'h313bab6d ;
    mem[8'h66] <= 32'hf923f82e ;
    mem[8'h67] <= 32'hbed436ef ;
    mem[8'h68] <= 32'h5bee0e79 ;
    mem[8'h69] <= 32'h1c19c0b8 ;
    mem[8'h6a] <= 32'hd40193fb ;
    mem[8'h6b] <= 32'h93f65d3a ;
    mem[8'h6c] <= 32'h40f028ca ;
    mem[8'h6d] <= 32'h707e60b ;
    mem[8'h6e] <= 32'hcf1fb548 ;
    mem[8'h6f] <= 32'h88e87b89 ;
    mem[8'h70] <= 32'h1aad9d3 ;
    mem[8'h71] <= 32'h465d1712 ;
    mem[8'h72] <= 32'h8e454451 ;
    mem[8'h73] <= 32'hc9b28a90 ;
    mem[8'h74] <= 32'h1ab4ff60 ;
    mem[8'h75] <= 32'h5d4331a1 ;
    mem[8'h76] <= 32'h955b62e2 ;
    mem[8'h77] <= 32'hd2acac23 ;
    mem[8'h78] <= 32'h379694b5 ;
    mem[8'h79] <= 32'h70615a74 ;
    mem[8'h7a] <= 32'hb8790937 ;
    mem[8'h7b] <= 32'hff8ec7f6 ;
    mem[8'h7c] <= 32'h2c88b206 ;
    mem[8'h7d] <= 32'h6b7f7cc7 ;
    mem[8'h7e] <= 32'ha3672f84 ;
    mem[8'h7f] <= 32'he490e145 ;
    mem[8'h80] <= 32'h6e87f0b9 ;
    mem[8'h81] <= 32'h29703e78 ;
    mem[8'h82] <= 32'he1686d3b ;
    mem[8'h83] <= 32'ha69fa3fa ;
    mem[8'h84] <= 32'h7599d60a ;
    mem[8'h85] <= 32'h326e18cb ;
    mem[8'h86] <= 32'hfa764b88 ;
    mem[8'h87] <= 32'hbd818549 ;
    mem[8'h88] <= 32'h58bbbddf ;
    mem[8'h89] <= 32'h1f4c731e ;
    mem[8'h8a] <= 32'hd754205d ;
    mem[8'h8b] <= 32'h90a3ee9c ;
    mem[8'h8c] <= 32'h43a59b6c ;
    mem[8'h8d] <= 32'h45255ad ;
    mem[8'h8e] <= 32'hcc4a06ee ;
    mem[8'h8f] <= 32'h8bbdc82f ;
    mem[8'h90] <= 32'h2ff6a75 ;
    mem[8'h91] <= 32'h4508a4b4 ;
    mem[8'h92] <= 32'h8d10f7f7 ;
    mem[8'h93] <= 32'hcae73936 ;
    mem[8'h94] <= 32'h19e14cc6 ;
    mem[8'h95] <= 32'h5e168207 ;
    mem[8'h96] <= 32'h960ed144 ;
    mem[8'h97] <= 32'hd1f91f85 ;
    mem[8'h98] <= 32'h34c32713 ;
    mem[8'h99] <= 32'h7334e9d2 ;
    mem[8'h9a] <= 32'hbb2cba91 ;
    mem[8'h9b] <= 32'hfcdb7450 ;
    mem[8'h9c] <= 32'h2fdd01a0 ;
    mem[8'h9d] <= 32'h682acf61 ;
    mem[8'h9e] <= 32'ha0329c22 ;
    mem[8'h9f] <= 32'he7c552e3 ;
    mem[8'ha0] <= 32'hb676c521 ;
    mem[8'ha1] <= 32'hf1810be0 ;
    mem[8'ha2] <= 32'h399958a3 ;
    mem[8'ha3] <= 32'h7e6e9662 ;
    mem[8'ha4] <= 32'had68e392 ;
    mem[8'ha5] <= 32'hea9f2d53 ;
    mem[8'ha6] <= 32'h22877e10 ;
    mem[8'ha7] <= 32'h6570b0d1 ;
    mem[8'ha8] <= 32'h804a8847 ;
    mem[8'ha9] <= 32'hc7bd4686 ;
    mem[8'haa] <= 32'hfa515c5 ;
    mem[8'hab] <= 32'h4852db04 ;
    mem[8'hac] <= 32'h9b54aef4 ;
    mem[8'had] <= 32'hdca36035 ;
    mem[8'hae] <= 32'h14bb3376 ;
    mem[8'haf] <= 32'h534cfdb7 ;
    mem[8'hb0] <= 32'hda0e5fed ;
    mem[8'hb1] <= 32'h9df9912c ;
    mem[8'hb2] <= 32'h55e1c26f ;
    mem[8'hb3] <= 32'h12160cae ;
    mem[8'hb4] <= 32'hc110795e ;
    mem[8'hb5] <= 32'h86e7b79f ;
    mem[8'hb6] <= 32'h4effe4dc ;
    mem[8'hb7] <= 32'h9082a1d ;
    mem[8'hb8] <= 32'hec32128b ;
    mem[8'hb9] <= 32'habc5dc4a ;
    mem[8'hba] <= 32'h63dd8f09 ;
    mem[8'hbb] <= 32'h242a41c8 ;
    mem[8'hbc] <= 32'hf72c3438 ;
    mem[8'hbd] <= 32'hb0dbfaf9 ;
    mem[8'hbe] <= 32'h78c3a9ba ;
    mem[8'hbf] <= 32'h3f34677b ;
    mem[8'hc0] <= 32'hdba4863e ;
    mem[8'hc1] <= 32'h9c5348ff ;
    mem[8'hc2] <= 32'h544b1bbc ;
    mem[8'hc3] <= 32'h13bcd57d ;
    mem[8'hc4] <= 32'hc0baa08d ;
    mem[8'hc5] <= 32'h874d6e4c ;
    mem[8'hc6] <= 32'h4f553d0f ;
    mem[8'hc7] <= 32'h8a2f3ce ;
    mem[8'hc8] <= 32'hed98cb58 ;
    mem[8'hc9] <= 32'haa6f0599 ;
    mem[8'hca] <= 32'h627756da ;
    mem[8'hcb] <= 32'h2580981b ;
    mem[8'hcc] <= 32'hf686edeb ;
    mem[8'hcd] <= 32'hb171232a ;
    mem[8'hce] <= 32'h79697069 ;
    mem[8'hcf] <= 32'h3e9ebea8 ;
    mem[8'hd0] <= 32'hb7dc1cf2 ;
    mem[8'hd1] <= 32'hf02bd233 ;
    mem[8'hd2] <= 32'h38338170 ;
    mem[8'hd3] <= 32'h7fc44fb1 ;
    mem[8'hd4] <= 32'hacc23a41 ;
    mem[8'hd5] <= 32'heb35f480 ;
    mem[8'hd6] <= 32'h232da7c3 ;
    mem[8'hd7] <= 32'h64da6902 ;
    mem[8'hd8] <= 32'h81e05194 ;
    mem[8'hd9] <= 32'hc6179f55 ;
    mem[8'hda] <= 32'he0fcc16 ;
    mem[8'hdb] <= 32'h49f802d7 ;
    mem[8'hdc] <= 32'h9afe7727 ;
    mem[8'hdd] <= 32'hdd09b9e6 ;
    mem[8'hde] <= 32'h1511eaa5 ;
    mem[8'hdf] <= 32'h52e62464 ;
    mem[8'he0] <= 32'h355b3a6 ;
    mem[8'he1] <= 32'h44a27d67 ;
    mem[8'he2] <= 32'h8cba2e24 ;
    mem[8'he3] <= 32'hcb4de0e5 ;
    mem[8'he4] <= 32'h184b9515 ;
    mem[8'he5] <= 32'h5fbc5bd4 ;
    mem[8'he6] <= 32'h97a40897 ;
    mem[8'he7] <= 32'hd053c656 ;
    mem[8'he8] <= 32'h3569fec0 ;
    mem[8'he9] <= 32'h729e3001 ;
    mem[8'hea] <= 32'hba866342 ;
    mem[8'heb] <= 32'hfd71ad83 ;
    mem[8'hec] <= 32'h2e77d873 ;
    mem[8'hed] <= 32'h698016b2 ;
    mem[8'hee] <= 32'ha19845f1 ;
    mem[8'hef] <= 32'he66f8b30 ;
    mem[8'hf0] <= 32'h6f2d296a ;
    mem[8'hf1] <= 32'h28dae7ab ;
    mem[8'hf2] <= 32'he0c2b4e8 ;
    mem[8'hf3] <= 32'ha7357a29 ;
    mem[8'hf4] <= 32'h74330fd9 ;
    mem[8'hf5] <= 32'h33c4c118 ;
    mem[8'hf6] <= 32'hfbdc925b ;
    mem[8'hf7] <= 32'hbc2b5c9a ;
    mem[8'hf8] <= 32'h5911640c ;
    mem[8'hf9] <= 32'h1ee6aacd ;
    mem[8'hfa] <= 32'hd6fef98e ;
    mem[8'hfb] <= 32'h9109374f ;
    mem[8'hfc] <= 32'h420f42bf ;
    mem[8'hfd] <= 32'h5f88c7e ;
    mem[8'hfe] <= 32'hcde0df3d ;
    mem[8'hff] <= 32'h8a1711fc ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
