module crctab_ev1
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'hd219c1dc ;
    mem[8'h2] <= 32'ha0f29e0f ;
    mem[8'h3] <= 32'h72eb5fd3 ;
    mem[8'h4] <= 32'h452421a9 ;
    mem[8'h5] <= 32'h973de075 ;
    mem[8'h6] <= 32'he5d6bfa6 ;
    mem[8'h7] <= 32'h37cf7e7a ;
    mem[8'h8] <= 32'h8a484352 ;
    mem[8'h9] <= 32'h5851828e ;
    mem[8'ha] <= 32'h2abadd5d ;
    mem[8'hb] <= 32'hf8a31c81 ;
    mem[8'hc] <= 32'hcf6c62fb ;
    mem[8'hd] <= 32'h1d75a327 ;
    mem[8'he] <= 32'h6f9efcf4 ;
    mem[8'hf] <= 32'hbd873d28 ;
    mem[8'h10] <= 32'h10519b13 ;
    mem[8'h11] <= 32'hc2485acf ;
    mem[8'h12] <= 32'hb0a3051c ;
    mem[8'h13] <= 32'h62bac4c0 ;
    mem[8'h14] <= 32'h5575baba ;
    mem[8'h15] <= 32'h876c7b66 ;
    mem[8'h16] <= 32'hf58724b5 ;
    mem[8'h17] <= 32'h279ee569 ;
    mem[8'h18] <= 32'h9a19d841 ;
    mem[8'h19] <= 32'h4800199d ;
    mem[8'h1a] <= 32'h3aeb464e ;
    mem[8'h1b] <= 32'he8f28792 ;
    mem[8'h1c] <= 32'hdf3df9e8 ;
    mem[8'h1d] <= 32'hd243834 ;
    mem[8'h1e] <= 32'h7fcf67e7 ;
    mem[8'h1f] <= 32'hadd6a63b ;
    mem[8'h20] <= 32'h20a33626 ;
    mem[8'h21] <= 32'hf2baf7fa ;
    mem[8'h22] <= 32'h8051a829 ;
    mem[8'h23] <= 32'h524869f5 ;
    mem[8'h24] <= 32'h6587178f ;
    mem[8'h25] <= 32'hb79ed653 ;
    mem[8'h26] <= 32'hc5758980 ;
    mem[8'h27] <= 32'h176c485c ;
    mem[8'h28] <= 32'haaeb7574 ;
    mem[8'h29] <= 32'h78f2b4a8 ;
    mem[8'h2a] <= 32'ha19eb7b ;
    mem[8'h2b] <= 32'hd8002aa7 ;
    mem[8'h2c] <= 32'hefcf54dd ;
    mem[8'h2d] <= 32'h3dd69501 ;
    mem[8'h2e] <= 32'h4f3dcad2 ;
    mem[8'h2f] <= 32'h9d240b0e ;
    mem[8'h30] <= 32'h30f2ad35 ;
    mem[8'h31] <= 32'he2eb6ce9 ;
    mem[8'h32] <= 32'h9000333a ;
    mem[8'h33] <= 32'h4219f2e6 ;
    mem[8'h34] <= 32'h75d68c9c ;
    mem[8'h35] <= 32'ha7cf4d40 ;
    mem[8'h36] <= 32'hd5241293 ;
    mem[8'h37] <= 32'h73dd34f ;
    mem[8'h38] <= 32'hbabaee67 ;
    mem[8'h39] <= 32'h68a32fbb ;
    mem[8'h3a] <= 32'h1a487068 ;
    mem[8'h3b] <= 32'hc851b1b4 ;
    mem[8'h3c] <= 32'hff9ecfce ;
    mem[8'h3d] <= 32'h2d870e12 ;
    mem[8'h3e] <= 32'h5f6c51c1 ;
    mem[8'h3f] <= 32'h8d75901d ;
    mem[8'h40] <= 32'h41466c4c ;
    mem[8'h41] <= 32'h935fad90 ;
    mem[8'h42] <= 32'he1b4f243 ;
    mem[8'h43] <= 32'h33ad339f ;
    mem[8'h44] <= 32'h4624de5 ;
    mem[8'h45] <= 32'hd67b8c39 ;
    mem[8'h46] <= 32'ha490d3ea ;
    mem[8'h47] <= 32'h76891236 ;
    mem[8'h48] <= 32'hcb0e2f1e ;
    mem[8'h49] <= 32'h1917eec2 ;
    mem[8'h4a] <= 32'h6bfcb111 ;
    mem[8'h4b] <= 32'hb9e570cd ;
    mem[8'h4c] <= 32'h8e2a0eb7 ;
    mem[8'h4d] <= 32'h5c33cf6b ;
    mem[8'h4e] <= 32'h2ed890b8 ;
    mem[8'h4f] <= 32'hfcc15164 ;
    mem[8'h50] <= 32'h5117f75f ;
    mem[8'h51] <= 32'h830e3683 ;
    mem[8'h52] <= 32'hf1e56950 ;
    mem[8'h53] <= 32'h23fca88c ;
    mem[8'h54] <= 32'h1433d6f6 ;
    mem[8'h55] <= 32'hc62a172a ;
    mem[8'h56] <= 32'hb4c148f9 ;
    mem[8'h57] <= 32'h66d88925 ;
    mem[8'h58] <= 32'hdb5fb40d ;
    mem[8'h59] <= 32'h94675d1 ;
    mem[8'h5a] <= 32'h7bad2a02 ;
    mem[8'h5b] <= 32'ha9b4ebde ;
    mem[8'h5c] <= 32'h9e7b95a4 ;
    mem[8'h5d] <= 32'h4c625478 ;
    mem[8'h5e] <= 32'h3e890bab ;
    mem[8'h5f] <= 32'hec90ca77 ;
    mem[8'h60] <= 32'h61e55a6a ;
    mem[8'h61] <= 32'hb3fc9bb6 ;
    mem[8'h62] <= 32'hc117c465 ;
    mem[8'h63] <= 32'h130e05b9 ;
    mem[8'h64] <= 32'h24c17bc3 ;
    mem[8'h65] <= 32'hf6d8ba1f ;
    mem[8'h66] <= 32'h8433e5cc ;
    mem[8'h67] <= 32'h562a2410 ;
    mem[8'h68] <= 32'hebad1938 ;
    mem[8'h69] <= 32'h39b4d8e4 ;
    mem[8'h6a] <= 32'h4b5f8737 ;
    mem[8'h6b] <= 32'h994646eb ;
    mem[8'h6c] <= 32'hae893891 ;
    mem[8'h6d] <= 32'h7c90f94d ;
    mem[8'h6e] <= 32'he7ba69e ;
    mem[8'h6f] <= 32'hdc626742 ;
    mem[8'h70] <= 32'h71b4c179 ;
    mem[8'h71] <= 32'ha3ad00a5 ;
    mem[8'h72] <= 32'hd1465f76 ;
    mem[8'h73] <= 32'h35f9eaa ;
    mem[8'h74] <= 32'h3490e0d0 ;
    mem[8'h75] <= 32'he689210c ;
    mem[8'h76] <= 32'h94627edf ;
    mem[8'h77] <= 32'h467bbf03 ;
    mem[8'h78] <= 32'hfbfc822b ;
    mem[8'h79] <= 32'h29e543f7 ;
    mem[8'h7a] <= 32'h5b0e1c24 ;
    mem[8'h7b] <= 32'h8917ddf8 ;
    mem[8'h7c] <= 32'hbed8a382 ;
    mem[8'h7d] <= 32'h6cc1625e ;
    mem[8'h7e] <= 32'h1e2a3d8d ;
    mem[8'h7f] <= 32'hcc33fc51 ;
    mem[8'h80] <= 32'h828cd898 ;
    mem[8'h81] <= 32'h50951944 ;
    mem[8'h82] <= 32'h227e4697 ;
    mem[8'h83] <= 32'hf067874b ;
    mem[8'h84] <= 32'hc7a8f931 ;
    mem[8'h85] <= 32'h15b138ed ;
    mem[8'h86] <= 32'h675a673e ;
    mem[8'h87] <= 32'hb543a6e2 ;
    mem[8'h88] <= 32'h8c49bca ;
    mem[8'h89] <= 32'hdadd5a16 ;
    mem[8'h8a] <= 32'ha83605c5 ;
    mem[8'h8b] <= 32'h7a2fc419 ;
    mem[8'h8c] <= 32'h4de0ba63 ;
    mem[8'h8d] <= 32'h9ff97bbf ;
    mem[8'h8e] <= 32'hed12246c ;
    mem[8'h8f] <= 32'h3f0be5b0 ;
    mem[8'h90] <= 32'h92dd438b ;
    mem[8'h91] <= 32'h40c48257 ;
    mem[8'h92] <= 32'h322fdd84 ;
    mem[8'h93] <= 32'he0361c58 ;
    mem[8'h94] <= 32'hd7f96222 ;
    mem[8'h95] <= 32'h5e0a3fe ;
    mem[8'h96] <= 32'h770bfc2d ;
    mem[8'h97] <= 32'ha5123df1 ;
    mem[8'h98] <= 32'h189500d9 ;
    mem[8'h99] <= 32'hca8cc105 ;
    mem[8'h9a] <= 32'hb8679ed6 ;
    mem[8'h9b] <= 32'h6a7e5f0a ;
    mem[8'h9c] <= 32'h5db12170 ;
    mem[8'h9d] <= 32'h8fa8e0ac ;
    mem[8'h9e] <= 32'hfd43bf7f ;
    mem[8'h9f] <= 32'h2f5a7ea3 ;
    mem[8'ha0] <= 32'ha22feebe ;
    mem[8'ha1] <= 32'h70362f62 ;
    mem[8'ha2] <= 32'h2dd70b1 ;
    mem[8'ha3] <= 32'hd0c4b16d ;
    mem[8'ha4] <= 32'he70bcf17 ;
    mem[8'ha5] <= 32'h35120ecb ;
    mem[8'ha6] <= 32'h47f95118 ;
    mem[8'ha7] <= 32'h95e090c4 ;
    mem[8'ha8] <= 32'h2867adec ;
    mem[8'ha9] <= 32'hfa7e6c30 ;
    mem[8'haa] <= 32'h889533e3 ;
    mem[8'hab] <= 32'h5a8cf23f ;
    mem[8'hac] <= 32'h6d438c45 ;
    mem[8'had] <= 32'hbf5a4d99 ;
    mem[8'hae] <= 32'hcdb1124a ;
    mem[8'haf] <= 32'h1fa8d396 ;
    mem[8'hb0] <= 32'hb27e75ad ;
    mem[8'hb1] <= 32'h6067b471 ;
    mem[8'hb2] <= 32'h128ceba2 ;
    mem[8'hb3] <= 32'hc0952a7e ;
    mem[8'hb4] <= 32'hf75a5404 ;
    mem[8'hb5] <= 32'h254395d8 ;
    mem[8'hb6] <= 32'h57a8ca0b ;
    mem[8'hb7] <= 32'h85b10bd7 ;
    mem[8'hb8] <= 32'h383636ff ;
    mem[8'hb9] <= 32'hea2ff723 ;
    mem[8'hba] <= 32'h98c4a8f0 ;
    mem[8'hbb] <= 32'h4add692c ;
    mem[8'hbc] <= 32'h7d121756 ;
    mem[8'hbd] <= 32'haf0bd68a ;
    mem[8'hbe] <= 32'hdde08959 ;
    mem[8'hbf] <= 32'hff94885 ;
    mem[8'hc0] <= 32'hc3cab4d4 ;
    mem[8'hc1] <= 32'h11d37508 ;
    mem[8'hc2] <= 32'h63382adb ;
    mem[8'hc3] <= 32'hb121eb07 ;
    mem[8'hc4] <= 32'h86ee957d ;
    mem[8'hc5] <= 32'h54f754a1 ;
    mem[8'hc6] <= 32'h261c0b72 ;
    mem[8'hc7] <= 32'hf405caae ;
    mem[8'hc8] <= 32'h4982f786 ;
    mem[8'hc9] <= 32'h9b9b365a ;
    mem[8'hca] <= 32'he9706989 ;
    mem[8'hcb] <= 32'h3b69a855 ;
    mem[8'hcc] <= 32'hca6d62f ;
    mem[8'hcd] <= 32'hdebf17f3 ;
    mem[8'hce] <= 32'hac544820 ;
    mem[8'hcf] <= 32'h7e4d89fc ;
    mem[8'hd0] <= 32'hd39b2fc7 ;
    mem[8'hd1] <= 32'h182ee1b ;
    mem[8'hd2] <= 32'h7369b1c8 ;
    mem[8'hd3] <= 32'ha1707014 ;
    mem[8'hd4] <= 32'h96bf0e6e ;
    mem[8'hd5] <= 32'h44a6cfb2 ;
    mem[8'hd6] <= 32'h364d9061 ;
    mem[8'hd7] <= 32'he45451bd ;
    mem[8'hd8] <= 32'h59d36c95 ;
    mem[8'hd9] <= 32'h8bcaad49 ;
    mem[8'hda] <= 32'hf921f29a ;
    mem[8'hdb] <= 32'h2b383346 ;
    mem[8'hdc] <= 32'h1cf74d3c ;
    mem[8'hdd] <= 32'hceee8ce0 ;
    mem[8'hde] <= 32'hbc05d333 ;
    mem[8'hdf] <= 32'h6e1c12ef ;
    mem[8'he0] <= 32'he36982f2 ;
    mem[8'he1] <= 32'h3170432e ;
    mem[8'he2] <= 32'h439b1cfd ;
    mem[8'he3] <= 32'h9182dd21 ;
    mem[8'he4] <= 32'ha64da35b ;
    mem[8'he5] <= 32'h74546287 ;
    mem[8'he6] <= 32'h6bf3d54 ;
    mem[8'he7] <= 32'hd4a6fc88 ;
    mem[8'he8] <= 32'h6921c1a0 ;
    mem[8'he9] <= 32'hbb38007c ;
    mem[8'hea] <= 32'hc9d35faf ;
    mem[8'heb] <= 32'h1bca9e73 ;
    mem[8'hec] <= 32'h2c05e009 ;
    mem[8'hed] <= 32'hfe1c21d5 ;
    mem[8'hee] <= 32'h8cf77e06 ;
    mem[8'hef] <= 32'h5eeebfda ;
    mem[8'hf0] <= 32'hf33819e1 ;
    mem[8'hf1] <= 32'h2121d83d ;
    mem[8'hf2] <= 32'h53ca87ee ;
    mem[8'hf3] <= 32'h81d34632 ;
    mem[8'hf4] <= 32'hb61c3848 ;
    mem[8'hf5] <= 32'h6405f994 ;
    mem[8'hf6] <= 32'h16eea647 ;
    mem[8'hf7] <= 32'hc4f7679b ;
    mem[8'hf8] <= 32'h79705ab3 ;
    mem[8'hf9] <= 32'hab699b6f ;
    mem[8'hfa] <= 32'hd982c4bc ;
    mem[8'hfb] <= 32'hb9b0560 ;
    mem[8'hfc] <= 32'h3c547b1a ;
    mem[8'hfd] <= 32'hee4dbac6 ;
    mem[8'hfe] <= 32'h9ca6e515 ;
    mem[8'hff] <= 32'h4ebf24c9 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
