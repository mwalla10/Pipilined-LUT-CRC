module crctab_ev7
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h5ba1dcca ;
    mem[8'h2] <= 32'hb743b994 ;
    mem[8'h3] <= 32'hece2655e ;
    mem[8'h4] <= 32'h6a466e9f ;
    mem[8'h5] <= 32'h31e7b255 ;
    mem[8'h6] <= 32'hdd05d70b ;
    mem[8'h7] <= 32'h86a40bc1 ;
    mem[8'h8] <= 32'hd48cdd3e ;
    mem[8'h9] <= 32'h8f2d01f4 ;
    mem[8'ha] <= 32'h63cf64aa ;
    mem[8'hb] <= 32'h386eb860 ;
    mem[8'hc] <= 32'hbecab3a1 ;
    mem[8'hd] <= 32'he56b6f6b ;
    mem[8'he] <= 32'h9890a35 ;
    mem[8'hf] <= 32'h5228d6ff ;
    mem[8'h10] <= 32'hadd8a7cb ;
    mem[8'h11] <= 32'hf6797b01 ;
    mem[8'h12] <= 32'h1a9b1e5f ;
    mem[8'h13] <= 32'h413ac295 ;
    mem[8'h14] <= 32'hc79ec954 ;
    mem[8'h15] <= 32'h9c3f159e ;
    mem[8'h16] <= 32'h70dd70c0 ;
    mem[8'h17] <= 32'h2b7cac0a ;
    mem[8'h18] <= 32'h79547af5 ;
    mem[8'h19] <= 32'h22f5a63f ;
    mem[8'h1a] <= 32'hce17c361 ;
    mem[8'h1b] <= 32'h95b61fab ;
    mem[8'h1c] <= 32'h1312146a ;
    mem[8'h1d] <= 32'h48b3c8a0 ;
    mem[8'h1e] <= 32'ha451adfe ;
    mem[8'h1f] <= 32'hfff07134 ;
    mem[8'h20] <= 32'h5f705221 ;
    mem[8'h21] <= 32'h4d18eeb ;
    mem[8'h22] <= 32'he833ebb5 ;
    mem[8'h23] <= 32'hb392377f ;
    mem[8'h24] <= 32'h35363cbe ;
    mem[8'h25] <= 32'h6e97e074 ;
    mem[8'h26] <= 32'h8275852a ;
    mem[8'h27] <= 32'hd9d459e0 ;
    mem[8'h28] <= 32'h8bfc8f1f ;
    mem[8'h29] <= 32'hd05d53d5 ;
    mem[8'h2a] <= 32'h3cbf368b ;
    mem[8'h2b] <= 32'h671eea41 ;
    mem[8'h2c] <= 32'he1bae180 ;
    mem[8'h2d] <= 32'hba1b3d4a ;
    mem[8'h2e] <= 32'h56f95814 ;
    mem[8'h2f] <= 32'hd5884de ;
    mem[8'h30] <= 32'hf2a8f5ea ;
    mem[8'h31] <= 32'ha9092920 ;
    mem[8'h32] <= 32'h45eb4c7e ;
    mem[8'h33] <= 32'h1e4a90b4 ;
    mem[8'h34] <= 32'h98ee9b75 ;
    mem[8'h35] <= 32'hc34f47bf ;
    mem[8'h36] <= 32'h2fad22e1 ;
    mem[8'h37] <= 32'h740cfe2b ;
    mem[8'h38] <= 32'h262428d4 ;
    mem[8'h39] <= 32'h7d85f41e ;
    mem[8'h3a] <= 32'h91679140 ;
    mem[8'h3b] <= 32'hcac64d8a ;
    mem[8'h3c] <= 32'h4c62464b ;
    mem[8'h3d] <= 32'h17c39a81 ;
    mem[8'h3e] <= 32'hfb21ffdf ;
    mem[8'h3f] <= 32'ha0802315 ;
    mem[8'h40] <= 32'hbee0a442 ;
    mem[8'h41] <= 32'he5417888 ;
    mem[8'h42] <= 32'h9a31dd6 ;
    mem[8'h43] <= 32'h5202c11c ;
    mem[8'h44] <= 32'hd4a6cadd ;
    mem[8'h45] <= 32'h8f071617 ;
    mem[8'h46] <= 32'h63e57349 ;
    mem[8'h47] <= 32'h3844af83 ;
    mem[8'h48] <= 32'h6a6c797c ;
    mem[8'h49] <= 32'h31cda5b6 ;
    mem[8'h4a] <= 32'hdd2fc0e8 ;
    mem[8'h4b] <= 32'h868e1c22 ;
    mem[8'h4c] <= 32'h2a17e3 ;
    mem[8'h4d] <= 32'h5b8bcb29 ;
    mem[8'h4e] <= 32'hb769ae77 ;
    mem[8'h4f] <= 32'hecc872bd ;
    mem[8'h50] <= 32'h13380389 ;
    mem[8'h51] <= 32'h4899df43 ;
    mem[8'h52] <= 32'ha47bba1d ;
    mem[8'h53] <= 32'hffda66d7 ;
    mem[8'h54] <= 32'h797e6d16 ;
    mem[8'h55] <= 32'h22dfb1dc ;
    mem[8'h56] <= 32'hce3dd482 ;
    mem[8'h57] <= 32'h959c0848 ;
    mem[8'h58] <= 32'hc7b4deb7 ;
    mem[8'h59] <= 32'h9c15027d ;
    mem[8'h5a] <= 32'h70f76723 ;
    mem[8'h5b] <= 32'h2b56bbe9 ;
    mem[8'h5c] <= 32'hadf2b028 ;
    mem[8'h5d] <= 32'hf6536ce2 ;
    mem[8'h5e] <= 32'h1ab109bc ;
    mem[8'h5f] <= 32'h4110d576 ;
    mem[8'h60] <= 32'he190f663 ;
    mem[8'h61] <= 32'hba312aa9 ;
    mem[8'h62] <= 32'h56d34ff7 ;
    mem[8'h63] <= 32'hd72933d ;
    mem[8'h64] <= 32'h8bd698fc ;
    mem[8'h65] <= 32'hd0774436 ;
    mem[8'h66] <= 32'h3c952168 ;
    mem[8'h67] <= 32'h6734fda2 ;
    mem[8'h68] <= 32'h351c2b5d ;
    mem[8'h69] <= 32'h6ebdf797 ;
    mem[8'h6a] <= 32'h825f92c9 ;
    mem[8'h6b] <= 32'hd9fe4e03 ;
    mem[8'h6c] <= 32'h5f5a45c2 ;
    mem[8'h6d] <= 32'h4fb9908 ;
    mem[8'h6e] <= 32'he819fc56 ;
    mem[8'h6f] <= 32'hb3b8209c ;
    mem[8'h70] <= 32'h4c4851a8 ;
    mem[8'h71] <= 32'h17e98d62 ;
    mem[8'h72] <= 32'hfb0be83c ;
    mem[8'h73] <= 32'ha0aa34f6 ;
    mem[8'h74] <= 32'h260e3f37 ;
    mem[8'h75] <= 32'h7dafe3fd ;
    mem[8'h76] <= 32'h914d86a3 ;
    mem[8'h77] <= 32'hcaec5a69 ;
    mem[8'h78] <= 32'h98c48c96 ;
    mem[8'h79] <= 32'hc365505c ;
    mem[8'h7a] <= 32'h2f873502 ;
    mem[8'h7b] <= 32'h7426e9c8 ;
    mem[8'h7c] <= 32'hf282e209 ;
    mem[8'h7d] <= 32'ha9233ec3 ;
    mem[8'h7e] <= 32'h45c15b9d ;
    mem[8'h7f] <= 32'h1e608757 ;
    mem[8'h80] <= 32'h79005533 ;
    mem[8'h81] <= 32'h22a189f9 ;
    mem[8'h82] <= 32'hce43eca7 ;
    mem[8'h83] <= 32'h95e2306d ;
    mem[8'h84] <= 32'h13463bac ;
    mem[8'h85] <= 32'h48e7e766 ;
    mem[8'h86] <= 32'ha4058238 ;
    mem[8'h87] <= 32'hffa45ef2 ;
    mem[8'h88] <= 32'had8c880d ;
    mem[8'h89] <= 32'hf62d54c7 ;
    mem[8'h8a] <= 32'h1acf3199 ;
    mem[8'h8b] <= 32'h416eed53 ;
    mem[8'h8c] <= 32'hc7cae692 ;
    mem[8'h8d] <= 32'h9c6b3a58 ;
    mem[8'h8e] <= 32'h70895f06 ;
    mem[8'h8f] <= 32'h2b2883cc ;
    mem[8'h90] <= 32'hd4d8f2f8 ;
    mem[8'h91] <= 32'h8f792e32 ;
    mem[8'h92] <= 32'h639b4b6c ;
    mem[8'h93] <= 32'h383a97a6 ;
    mem[8'h94] <= 32'hbe9e9c67 ;
    mem[8'h95] <= 32'he53f40ad ;
    mem[8'h96] <= 32'h9dd25f3 ;
    mem[8'h97] <= 32'h527cf939 ;
    mem[8'h98] <= 32'h542fc6 ;
    mem[8'h99] <= 32'h5bf5f30c ;
    mem[8'h9a] <= 32'hb7179652 ;
    mem[8'h9b] <= 32'hecb64a98 ;
    mem[8'h9c] <= 32'h6a124159 ;
    mem[8'h9d] <= 32'h31b39d93 ;
    mem[8'h9e] <= 32'hdd51f8cd ;
    mem[8'h9f] <= 32'h86f02407 ;
    mem[8'ha0] <= 32'h26700712 ;
    mem[8'ha1] <= 32'h7dd1dbd8 ;
    mem[8'ha2] <= 32'h9133be86 ;
    mem[8'ha3] <= 32'hca92624c ;
    mem[8'ha4] <= 32'h4c36698d ;
    mem[8'ha5] <= 32'h1797b547 ;
    mem[8'ha6] <= 32'hfb75d019 ;
    mem[8'ha7] <= 32'ha0d40cd3 ;
    mem[8'ha8] <= 32'hf2fcda2c ;
    mem[8'ha9] <= 32'ha95d06e6 ;
    mem[8'haa] <= 32'h45bf63b8 ;
    mem[8'hab] <= 32'h1e1ebf72 ;
    mem[8'hac] <= 32'h98bab4b3 ;
    mem[8'had] <= 32'hc31b6879 ;
    mem[8'hae] <= 32'h2ff90d27 ;
    mem[8'haf] <= 32'h7458d1ed ;
    mem[8'hb0] <= 32'h8ba8a0d9 ;
    mem[8'hb1] <= 32'hd0097c13 ;
    mem[8'hb2] <= 32'h3ceb194d ;
    mem[8'hb3] <= 32'h674ac587 ;
    mem[8'hb4] <= 32'he1eece46 ;
    mem[8'hb5] <= 32'hba4f128c ;
    mem[8'hb6] <= 32'h56ad77d2 ;
    mem[8'hb7] <= 32'hd0cab18 ;
    mem[8'hb8] <= 32'h5f247de7 ;
    mem[8'hb9] <= 32'h485a12d ;
    mem[8'hba] <= 32'he867c473 ;
    mem[8'hbb] <= 32'hb3c618b9 ;
    mem[8'hbc] <= 32'h35621378 ;
    mem[8'hbd] <= 32'h6ec3cfb2 ;
    mem[8'hbe] <= 32'h8221aaec ;
    mem[8'hbf] <= 32'hd9807626 ;
    mem[8'hc0] <= 32'hc7e0f171 ;
    mem[8'hc1] <= 32'h9c412dbb ;
    mem[8'hc2] <= 32'h70a348e5 ;
    mem[8'hc3] <= 32'h2b02942f ;
    mem[8'hc4] <= 32'hada69fee ;
    mem[8'hc5] <= 32'hf6074324 ;
    mem[8'hc6] <= 32'h1ae5267a ;
    mem[8'hc7] <= 32'h4144fab0 ;
    mem[8'hc8] <= 32'h136c2c4f ;
    mem[8'hc9] <= 32'h48cdf085 ;
    mem[8'hca] <= 32'ha42f95db ;
    mem[8'hcb] <= 32'hff8e4911 ;
    mem[8'hcc] <= 32'h792a42d0 ;
    mem[8'hcd] <= 32'h228b9e1a ;
    mem[8'hce] <= 32'hce69fb44 ;
    mem[8'hcf] <= 32'h95c8278e ;
    mem[8'hd0] <= 32'h6a3856ba ;
    mem[8'hd1] <= 32'h31998a70 ;
    mem[8'hd2] <= 32'hdd7bef2e ;
    mem[8'hd3] <= 32'h86da33e4 ;
    mem[8'hd4] <= 32'h7e3825 ;
    mem[8'hd5] <= 32'h5bdfe4ef ;
    mem[8'hd6] <= 32'hb73d81b1 ;
    mem[8'hd7] <= 32'hec9c5d7b ;
    mem[8'hd8] <= 32'hbeb48b84 ;
    mem[8'hd9] <= 32'he515574e ;
    mem[8'hda] <= 32'h9f73210 ;
    mem[8'hdb] <= 32'h5256eeda ;
    mem[8'hdc] <= 32'hd4f2e51b ;
    mem[8'hdd] <= 32'h8f5339d1 ;
    mem[8'hde] <= 32'h63b15c8f ;
    mem[8'hdf] <= 32'h38108045 ;
    mem[8'he0] <= 32'h9890a350 ;
    mem[8'he1] <= 32'hc3317f9a ;
    mem[8'he2] <= 32'h2fd31ac4 ;
    mem[8'he3] <= 32'h7472c60e ;
    mem[8'he4] <= 32'hf2d6cdcf ;
    mem[8'he5] <= 32'ha9771105 ;
    mem[8'he6] <= 32'h4595745b ;
    mem[8'he7] <= 32'h1e34a891 ;
    mem[8'he8] <= 32'h4c1c7e6e ;
    mem[8'he9] <= 32'h17bda2a4 ;
    mem[8'hea] <= 32'hfb5fc7fa ;
    mem[8'heb] <= 32'ha0fe1b30 ;
    mem[8'hec] <= 32'h265a10f1 ;
    mem[8'hed] <= 32'h7dfbcc3b ;
    mem[8'hee] <= 32'h9119a965 ;
    mem[8'hef] <= 32'hcab875af ;
    mem[8'hf0] <= 32'h3548049b ;
    mem[8'hf1] <= 32'h6ee9d851 ;
    mem[8'hf2] <= 32'h820bbd0f ;
    mem[8'hf3] <= 32'hd9aa61c5 ;
    mem[8'hf4] <= 32'h5f0e6a04 ;
    mem[8'hf5] <= 32'h4afb6ce ;
    mem[8'hf6] <= 32'he84dd390 ;
    mem[8'hf7] <= 32'hb3ec0f5a ;
    mem[8'hf8] <= 32'he1c4d9a5 ;
    mem[8'hf9] <= 32'hba65056f ;
    mem[8'hfa] <= 32'h56876031 ;
    mem[8'hfb] <= 32'hd26bcfb ;
    mem[8'hfc] <= 32'h8b82b73a ;
    mem[8'hfd] <= 32'hd0236bf0 ;
    mem[8'hfe] <= 32'h3cc10eae ;
    mem[8'hff] <= 32'h6760d264 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
