module crctab_ev30
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h218e0c78 ;
    mem[8'h2] <= 32'h431c18f0 ;
    mem[8'h3] <= 32'h62921488 ;
    mem[8'h4] <= 32'h863831e0 ;
    mem[8'h5] <= 32'ha7b63d98 ;
    mem[8'h6] <= 32'hc5242910 ;
    mem[8'h7] <= 32'he4aa2568 ;
    mem[8'h8] <= 32'h8b17e77 ;
    mem[8'h9] <= 32'h293f720f ;
    mem[8'ha] <= 32'h4bad6687 ;
    mem[8'hb] <= 32'h6a236aff ;
    mem[8'hc] <= 32'h8e894f97 ;
    mem[8'hd] <= 32'haf0743ef ;
    mem[8'he] <= 32'hcd955767 ;
    mem[8'hf] <= 32'hec1b5b1f ;
    mem[8'h10] <= 32'h1162fcee ;
    mem[8'h11] <= 32'h30ecf096 ;
    mem[8'h12] <= 32'h527ee41e ;
    mem[8'h13] <= 32'h73f0e866 ;
    mem[8'h14] <= 32'h975acd0e ;
    mem[8'h15] <= 32'hb6d4c176 ;
    mem[8'h16] <= 32'hd446d5fe ;
    mem[8'h17] <= 32'hf5c8d986 ;
    mem[8'h18] <= 32'h19d38299 ;
    mem[8'h19] <= 32'h385d8ee1 ;
    mem[8'h1a] <= 32'h5acf9a69 ;
    mem[8'h1b] <= 32'h7b419611 ;
    mem[8'h1c] <= 32'h9febb379 ;
    mem[8'h1d] <= 32'hbe65bf01 ;
    mem[8'h1e] <= 32'hdcf7ab89 ;
    mem[8'h1f] <= 32'hfd79a7f1 ;
    mem[8'h20] <= 32'h22c5f9dc ;
    mem[8'h21] <= 32'h34bf5a4 ;
    mem[8'h22] <= 32'h61d9e12c ;
    mem[8'h23] <= 32'h4057ed54 ;
    mem[8'h24] <= 32'ha4fdc83c ;
    mem[8'h25] <= 32'h8573c444 ;
    mem[8'h26] <= 32'he7e1d0cc ;
    mem[8'h27] <= 32'hc66fdcb4 ;
    mem[8'h28] <= 32'h2a7487ab ;
    mem[8'h29] <= 32'hbfa8bd3 ;
    mem[8'h2a] <= 32'h69689f5b ;
    mem[8'h2b] <= 32'h48e69323 ;
    mem[8'h2c] <= 32'hac4cb64b ;
    mem[8'h2d] <= 32'h8dc2ba33 ;
    mem[8'h2e] <= 32'hef50aebb ;
    mem[8'h2f] <= 32'hcedea2c3 ;
    mem[8'h30] <= 32'h33a70532 ;
    mem[8'h31] <= 32'h1229094a ;
    mem[8'h32] <= 32'h70bb1dc2 ;
    mem[8'h33] <= 32'h513511ba ;
    mem[8'h34] <= 32'hb59f34d2 ;
    mem[8'h35] <= 32'h941138aa ;
    mem[8'h36] <= 32'hf6832c22 ;
    mem[8'h37] <= 32'hd70d205a ;
    mem[8'h38] <= 32'h3b167b45 ;
    mem[8'h39] <= 32'h1a98773d ;
    mem[8'h3a] <= 32'h780a63b5 ;
    mem[8'h3b] <= 32'h59846fcd ;
    mem[8'h3c] <= 32'hbd2e4aa5 ;
    mem[8'h3d] <= 32'h9ca046dd ;
    mem[8'h3e] <= 32'hfe325255 ;
    mem[8'h3f] <= 32'hdfbc5e2d ;
    mem[8'h40] <= 32'h458bf3b8 ;
    mem[8'h41] <= 32'h6405ffc0 ;
    mem[8'h42] <= 32'h697eb48 ;
    mem[8'h43] <= 32'h2719e730 ;
    mem[8'h44] <= 32'hc3b3c258 ;
    mem[8'h45] <= 32'he23dce20 ;
    mem[8'h46] <= 32'h80afdaa8 ;
    mem[8'h47] <= 32'ha121d6d0 ;
    mem[8'h48] <= 32'h4d3a8dcf ;
    mem[8'h49] <= 32'h6cb481b7 ;
    mem[8'h4a] <= 32'he26953f ;
    mem[8'h4b] <= 32'h2fa89947 ;
    mem[8'h4c] <= 32'hcb02bc2f ;
    mem[8'h4d] <= 32'hea8cb057 ;
    mem[8'h4e] <= 32'h881ea4df ;
    mem[8'h4f] <= 32'ha990a8a7 ;
    mem[8'h50] <= 32'h54e90f56 ;
    mem[8'h51] <= 32'h7567032e ;
    mem[8'h52] <= 32'h17f517a6 ;
    mem[8'h53] <= 32'h367b1bde ;
    mem[8'h54] <= 32'hd2d13eb6 ;
    mem[8'h55] <= 32'hf35f32ce ;
    mem[8'h56] <= 32'h91cd2646 ;
    mem[8'h57] <= 32'hb0432a3e ;
    mem[8'h58] <= 32'h5c587121 ;
    mem[8'h59] <= 32'h7dd67d59 ;
    mem[8'h5a] <= 32'h1f4469d1 ;
    mem[8'h5b] <= 32'h3eca65a9 ;
    mem[8'h5c] <= 32'hda6040c1 ;
    mem[8'h5d] <= 32'hfbee4cb9 ;
    mem[8'h5e] <= 32'h997c5831 ;
    mem[8'h5f] <= 32'hb8f25449 ;
    mem[8'h60] <= 32'h674e0a64 ;
    mem[8'h61] <= 32'h46c0061c ;
    mem[8'h62] <= 32'h24521294 ;
    mem[8'h63] <= 32'h5dc1eec ;
    mem[8'h64] <= 32'he1763b84 ;
    mem[8'h65] <= 32'hc0f837fc ;
    mem[8'h66] <= 32'ha26a2374 ;
    mem[8'h67] <= 32'h83e42f0c ;
    mem[8'h68] <= 32'h6fff7413 ;
    mem[8'h69] <= 32'h4e71786b ;
    mem[8'h6a] <= 32'h2ce36ce3 ;
    mem[8'h6b] <= 32'hd6d609b ;
    mem[8'h6c] <= 32'he9c745f3 ;
    mem[8'h6d] <= 32'hc849498b ;
    mem[8'h6e] <= 32'haadb5d03 ;
    mem[8'h6f] <= 32'h8b55517b ;
    mem[8'h70] <= 32'h762cf68a ;
    mem[8'h71] <= 32'h57a2faf2 ;
    mem[8'h72] <= 32'h3530ee7a ;
    mem[8'h73] <= 32'h14bee202 ;
    mem[8'h74] <= 32'hf014c76a ;
    mem[8'h75] <= 32'hd19acb12 ;
    mem[8'h76] <= 32'hb308df9a ;
    mem[8'h77] <= 32'h9286d3e2 ;
    mem[8'h78] <= 32'h7e9d88fd ;
    mem[8'h79] <= 32'h5f138485 ;
    mem[8'h7a] <= 32'h3d81900d ;
    mem[8'h7b] <= 32'h1c0f9c75 ;
    mem[8'h7c] <= 32'hf8a5b91d ;
    mem[8'h7d] <= 32'hd92bb565 ;
    mem[8'h7e] <= 32'hbbb9a1ed ;
    mem[8'h7f] <= 32'h9a37ad95 ;
    mem[8'h80] <= 32'h8b17e770 ;
    mem[8'h81] <= 32'haa99eb08 ;
    mem[8'h82] <= 32'hc80bff80 ;
    mem[8'h83] <= 32'he985f3f8 ;
    mem[8'h84] <= 32'hd2fd690 ;
    mem[8'h85] <= 32'h2ca1dae8 ;
    mem[8'h86] <= 32'h4e33ce60 ;
    mem[8'h87] <= 32'h6fbdc218 ;
    mem[8'h88] <= 32'h83a69907 ;
    mem[8'h89] <= 32'ha228957f ;
    mem[8'h8a] <= 32'hc0ba81f7 ;
    mem[8'h8b] <= 32'he1348d8f ;
    mem[8'h8c] <= 32'h59ea8e7 ;
    mem[8'h8d] <= 32'h2410a49f ;
    mem[8'h8e] <= 32'h4682b017 ;
    mem[8'h8f] <= 32'h670cbc6f ;
    mem[8'h90] <= 32'h9a751b9e ;
    mem[8'h91] <= 32'hbbfb17e6 ;
    mem[8'h92] <= 32'hd969036e ;
    mem[8'h93] <= 32'hf8e70f16 ;
    mem[8'h94] <= 32'h1c4d2a7e ;
    mem[8'h95] <= 32'h3dc32606 ;
    mem[8'h96] <= 32'h5f51328e ;
    mem[8'h97] <= 32'h7edf3ef6 ;
    mem[8'h98] <= 32'h92c465e9 ;
    mem[8'h99] <= 32'hb34a6991 ;
    mem[8'h9a] <= 32'hd1d87d19 ;
    mem[8'h9b] <= 32'hf0567161 ;
    mem[8'h9c] <= 32'h14fc5409 ;
    mem[8'h9d] <= 32'h35725871 ;
    mem[8'h9e] <= 32'h57e04cf9 ;
    mem[8'h9f] <= 32'h766e4081 ;
    mem[8'ha0] <= 32'ha9d21eac ;
    mem[8'ha1] <= 32'h885c12d4 ;
    mem[8'ha2] <= 32'heace065c ;
    mem[8'ha3] <= 32'hcb400a24 ;
    mem[8'ha4] <= 32'h2fea2f4c ;
    mem[8'ha5] <= 32'he642334 ;
    mem[8'ha6] <= 32'h6cf637bc ;
    mem[8'ha7] <= 32'h4d783bc4 ;
    mem[8'ha8] <= 32'ha16360db ;
    mem[8'ha9] <= 32'h80ed6ca3 ;
    mem[8'haa] <= 32'he27f782b ;
    mem[8'hab] <= 32'hc3f17453 ;
    mem[8'hac] <= 32'h275b513b ;
    mem[8'had] <= 32'h6d55d43 ;
    mem[8'hae] <= 32'h644749cb ;
    mem[8'haf] <= 32'h45c945b3 ;
    mem[8'hb0] <= 32'hb8b0e242 ;
    mem[8'hb1] <= 32'h993eee3a ;
    mem[8'hb2] <= 32'hfbacfab2 ;
    mem[8'hb3] <= 32'hda22f6ca ;
    mem[8'hb4] <= 32'h3e88d3a2 ;
    mem[8'hb5] <= 32'h1f06dfda ;
    mem[8'hb6] <= 32'h7d94cb52 ;
    mem[8'hb7] <= 32'h5c1ac72a ;
    mem[8'hb8] <= 32'hb0019c35 ;
    mem[8'hb9] <= 32'h918f904d ;
    mem[8'hba] <= 32'hf31d84c5 ;
    mem[8'hbb] <= 32'hd29388bd ;
    mem[8'hbc] <= 32'h3639add5 ;
    mem[8'hbd] <= 32'h17b7a1ad ;
    mem[8'hbe] <= 32'h7525b525 ;
    mem[8'hbf] <= 32'h54abb95d ;
    mem[8'hc0] <= 32'hce9c14c8 ;
    mem[8'hc1] <= 32'hef1218b0 ;
    mem[8'hc2] <= 32'h8d800c38 ;
    mem[8'hc3] <= 32'hac0e0040 ;
    mem[8'hc4] <= 32'h48a42528 ;
    mem[8'hc5] <= 32'h692a2950 ;
    mem[8'hc6] <= 32'hbb83dd8 ;
    mem[8'hc7] <= 32'h2a3631a0 ;
    mem[8'hc8] <= 32'hc62d6abf ;
    mem[8'hc9] <= 32'he7a366c7 ;
    mem[8'hca] <= 32'h8531724f ;
    mem[8'hcb] <= 32'ha4bf7e37 ;
    mem[8'hcc] <= 32'h40155b5f ;
    mem[8'hcd] <= 32'h619b5727 ;
    mem[8'hce] <= 32'h30943af ;
    mem[8'hcf] <= 32'h22874fd7 ;
    mem[8'hd0] <= 32'hdffee826 ;
    mem[8'hd1] <= 32'hfe70e45e ;
    mem[8'hd2] <= 32'h9ce2f0d6 ;
    mem[8'hd3] <= 32'hbd6cfcae ;
    mem[8'hd4] <= 32'h59c6d9c6 ;
    mem[8'hd5] <= 32'h7848d5be ;
    mem[8'hd6] <= 32'h1adac136 ;
    mem[8'hd7] <= 32'h3b54cd4e ;
    mem[8'hd8] <= 32'hd74f9651 ;
    mem[8'hd9] <= 32'hf6c19a29 ;
    mem[8'hda] <= 32'h94538ea1 ;
    mem[8'hdb] <= 32'hb5dd82d9 ;
    mem[8'hdc] <= 32'h5177a7b1 ;
    mem[8'hdd] <= 32'h70f9abc9 ;
    mem[8'hde] <= 32'h126bbf41 ;
    mem[8'hdf] <= 32'h33e5b339 ;
    mem[8'he0] <= 32'hec59ed14 ;
    mem[8'he1] <= 32'hcdd7e16c ;
    mem[8'he2] <= 32'haf45f5e4 ;
    mem[8'he3] <= 32'h8ecbf99c ;
    mem[8'he4] <= 32'h6a61dcf4 ;
    mem[8'he5] <= 32'h4befd08c ;
    mem[8'he6] <= 32'h297dc404 ;
    mem[8'he7] <= 32'h8f3c87c ;
    mem[8'he8] <= 32'he4e89363 ;
    mem[8'he9] <= 32'hc5669f1b ;
    mem[8'hea] <= 32'ha7f48b93 ;
    mem[8'heb] <= 32'h867a87eb ;
    mem[8'hec] <= 32'h62d0a283 ;
    mem[8'hed] <= 32'h435eaefb ;
    mem[8'hee] <= 32'h21ccba73 ;
    mem[8'hef] <= 32'h42b60b ;
    mem[8'hf0] <= 32'hfd3b11fa ;
    mem[8'hf1] <= 32'hdcb51d82 ;
    mem[8'hf2] <= 32'hbe27090a ;
    mem[8'hf3] <= 32'h9fa90572 ;
    mem[8'hf4] <= 32'h7b03201a ;
    mem[8'hf5] <= 32'h5a8d2c62 ;
    mem[8'hf6] <= 32'h381f38ea ;
    mem[8'hf7] <= 32'h19913492 ;
    mem[8'hf8] <= 32'hf58a6f8d ;
    mem[8'hf9] <= 32'hd40463f5 ;
    mem[8'hfa] <= 32'hb696777d ;
    mem[8'hfb] <= 32'h97187b05 ;
    mem[8'hfc] <= 32'h73b25e6d ;
    mem[8'hfd] <= 32'h523c5215 ;
    mem[8'hfe] <= 32'h30ae469d ;
    mem[8'hff] <= 32'h11204ae5 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
