module crctab_ev22
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h64c29d0 ;
    mem[8'h2] <= 32'hc9853a0 ;
    mem[8'h3] <= 32'had47a70 ;
    mem[8'h4] <= 32'h1930a740 ;
    mem[8'h5] <= 32'h1f7c8e90 ;
    mem[8'h6] <= 32'h15a8f4e0 ;
    mem[8'h7] <= 32'h13e4dd30 ;
    mem[8'h8] <= 32'h32614e80 ;
    mem[8'h9] <= 32'h342d6750 ;
    mem[8'ha] <= 32'h3ef91d20 ;
    mem[8'hb] <= 32'h38b534f0 ;
    mem[8'hc] <= 32'h2b51e9c0 ;
    mem[8'hd] <= 32'h2d1dc010 ;
    mem[8'he] <= 32'h27c9ba60 ;
    mem[8'hf] <= 32'h218593b0 ;
    mem[8'h10] <= 32'h64c29d00 ;
    mem[8'h11] <= 32'h628eb4d0 ;
    mem[8'h12] <= 32'h685acea0 ;
    mem[8'h13] <= 32'h6e16e770 ;
    mem[8'h14] <= 32'h7df23a40 ;
    mem[8'h15] <= 32'h7bbe1390 ;
    mem[8'h16] <= 32'h716a69e0 ;
    mem[8'h17] <= 32'h77264030 ;
    mem[8'h18] <= 32'h56a3d380 ;
    mem[8'h19] <= 32'h50effa50 ;
    mem[8'h1a] <= 32'h5a3b8020 ;
    mem[8'h1b] <= 32'h5c77a9f0 ;
    mem[8'h1c] <= 32'h4f9374c0 ;
    mem[8'h1d] <= 32'h49df5d10 ;
    mem[8'h1e] <= 32'h430b2760 ;
    mem[8'h1f] <= 32'h45470eb0 ;
    mem[8'h20] <= 32'hc9853a00 ;
    mem[8'h21] <= 32'hcfc913d0 ;
    mem[8'h22] <= 32'hc51d69a0 ;
    mem[8'h23] <= 32'hc3514070 ;
    mem[8'h24] <= 32'hd0b59d40 ;
    mem[8'h25] <= 32'hd6f9b490 ;
    mem[8'h26] <= 32'hdc2dcee0 ;
    mem[8'h27] <= 32'hda61e730 ;
    mem[8'h28] <= 32'hfbe47480 ;
    mem[8'h29] <= 32'hfda85d50 ;
    mem[8'h2a] <= 32'hf77c2720 ;
    mem[8'h2b] <= 32'hf1300ef0 ;
    mem[8'h2c] <= 32'he2d4d3c0 ;
    mem[8'h2d] <= 32'he498fa10 ;
    mem[8'h2e] <= 32'hee4c8060 ;
    mem[8'h2f] <= 32'he800a9b0 ;
    mem[8'h30] <= 32'had47a700 ;
    mem[8'h31] <= 32'hab0b8ed0 ;
    mem[8'h32] <= 32'ha1dff4a0 ;
    mem[8'h33] <= 32'ha793dd70 ;
    mem[8'h34] <= 32'hb4770040 ;
    mem[8'h35] <= 32'hb23b2990 ;
    mem[8'h36] <= 32'hb8ef53e0 ;
    mem[8'h37] <= 32'hbea37a30 ;
    mem[8'h38] <= 32'h9f26e980 ;
    mem[8'h39] <= 32'h996ac050 ;
    mem[8'h3a] <= 32'h93beba20 ;
    mem[8'h3b] <= 32'h95f293f0 ;
    mem[8'h3c] <= 32'h86164ec0 ;
    mem[8'h3d] <= 32'h805a6710 ;
    mem[8'h3e] <= 32'h8a8e1d60 ;
    mem[8'h3f] <= 32'h8cc234b0 ;
    mem[8'h40] <= 32'h97cb69b7 ;
    mem[8'h41] <= 32'h91874067 ;
    mem[8'h42] <= 32'h9b533a17 ;
    mem[8'h43] <= 32'h9d1f13c7 ;
    mem[8'h44] <= 32'h8efbcef7 ;
    mem[8'h45] <= 32'h88b7e727 ;
    mem[8'h46] <= 32'h82639d57 ;
    mem[8'h47] <= 32'h842fb487 ;
    mem[8'h48] <= 32'ha5aa2737 ;
    mem[8'h49] <= 32'ha3e60ee7 ;
    mem[8'h4a] <= 32'ha9327497 ;
    mem[8'h4b] <= 32'haf7e5d47 ;
    mem[8'h4c] <= 32'hbc9a8077 ;
    mem[8'h4d] <= 32'hbad6a9a7 ;
    mem[8'h4e] <= 32'hb002d3d7 ;
    mem[8'h4f] <= 32'hb64efa07 ;
    mem[8'h50] <= 32'hf309f4b7 ;
    mem[8'h51] <= 32'hf545dd67 ;
    mem[8'h52] <= 32'hff91a717 ;
    mem[8'h53] <= 32'hf9dd8ec7 ;
    mem[8'h54] <= 32'hea3953f7 ;
    mem[8'h55] <= 32'hec757a27 ;
    mem[8'h56] <= 32'he6a10057 ;
    mem[8'h57] <= 32'he0ed2987 ;
    mem[8'h58] <= 32'hc168ba37 ;
    mem[8'h59] <= 32'hc72493e7 ;
    mem[8'h5a] <= 32'hcdf0e997 ;
    mem[8'h5b] <= 32'hcbbcc047 ;
    mem[8'h5c] <= 32'hd8581d77 ;
    mem[8'h5d] <= 32'hde1434a7 ;
    mem[8'h5e] <= 32'hd4c04ed7 ;
    mem[8'h5f] <= 32'hd28c6707 ;
    mem[8'h60] <= 32'h5e4e53b7 ;
    mem[8'h61] <= 32'h58027a67 ;
    mem[8'h62] <= 32'h52d60017 ;
    mem[8'h63] <= 32'h549a29c7 ;
    mem[8'h64] <= 32'h477ef4f7 ;
    mem[8'h65] <= 32'h4132dd27 ;
    mem[8'h66] <= 32'h4be6a757 ;
    mem[8'h67] <= 32'h4daa8e87 ;
    mem[8'h68] <= 32'h6c2f1d37 ;
    mem[8'h69] <= 32'h6a6334e7 ;
    mem[8'h6a] <= 32'h60b74e97 ;
    mem[8'h6b] <= 32'h66fb6747 ;
    mem[8'h6c] <= 32'h751fba77 ;
    mem[8'h6d] <= 32'h735393a7 ;
    mem[8'h6e] <= 32'h7987e9d7 ;
    mem[8'h6f] <= 32'h7fcbc007 ;
    mem[8'h70] <= 32'h3a8cceb7 ;
    mem[8'h71] <= 32'h3cc0e767 ;
    mem[8'h72] <= 32'h36149d17 ;
    mem[8'h73] <= 32'h3058b4c7 ;
    mem[8'h74] <= 32'h23bc69f7 ;
    mem[8'h75] <= 32'h25f04027 ;
    mem[8'h76] <= 32'h2f243a57 ;
    mem[8'h77] <= 32'h29681387 ;
    mem[8'h78] <= 32'h8ed8037 ;
    mem[8'h79] <= 32'hea1a9e7 ;
    mem[8'h7a] <= 32'h475d397 ;
    mem[8'h7b] <= 32'h239fa47 ;
    mem[8'h7c] <= 32'h11dd2777 ;
    mem[8'h7d] <= 32'h17910ea7 ;
    mem[8'h7e] <= 32'h1d4574d7 ;
    mem[8'h7f] <= 32'h1b095d07 ;
    mem[8'h80] <= 32'h2b57ced9 ;
    mem[8'h81] <= 32'h2d1be709 ;
    mem[8'h82] <= 32'h27cf9d79 ;
    mem[8'h83] <= 32'h2183b4a9 ;
    mem[8'h84] <= 32'h32676999 ;
    mem[8'h85] <= 32'h342b4049 ;
    mem[8'h86] <= 32'h3eff3a39 ;
    mem[8'h87] <= 32'h38b313e9 ;
    mem[8'h88] <= 32'h19368059 ;
    mem[8'h89] <= 32'h1f7aa989 ;
    mem[8'h8a] <= 32'h15aed3f9 ;
    mem[8'h8b] <= 32'h13e2fa29 ;
    mem[8'h8c] <= 32'h62719 ;
    mem[8'h8d] <= 32'h64a0ec9 ;
    mem[8'h8e] <= 32'hc9e74b9 ;
    mem[8'h8f] <= 32'had25d69 ;
    mem[8'h90] <= 32'h4f9553d9 ;
    mem[8'h91] <= 32'h49d97a09 ;
    mem[8'h92] <= 32'h430d0079 ;
    mem[8'h93] <= 32'h454129a9 ;
    mem[8'h94] <= 32'h56a5f499 ;
    mem[8'h95] <= 32'h50e9dd49 ;
    mem[8'h96] <= 32'h5a3da739 ;
    mem[8'h97] <= 32'h5c718ee9 ;
    mem[8'h98] <= 32'h7df41d59 ;
    mem[8'h99] <= 32'h7bb83489 ;
    mem[8'h9a] <= 32'h716c4ef9 ;
    mem[8'h9b] <= 32'h77206729 ;
    mem[8'h9c] <= 32'h64c4ba19 ;
    mem[8'h9d] <= 32'h628893c9 ;
    mem[8'h9e] <= 32'h685ce9b9 ;
    mem[8'h9f] <= 32'h6e10c069 ;
    mem[8'ha0] <= 32'he2d2f4d9 ;
    mem[8'ha1] <= 32'he49edd09 ;
    mem[8'ha2] <= 32'hee4aa779 ;
    mem[8'ha3] <= 32'he8068ea9 ;
    mem[8'ha4] <= 32'hfbe25399 ;
    mem[8'ha5] <= 32'hfdae7a49 ;
    mem[8'ha6] <= 32'hf77a0039 ;
    mem[8'ha7] <= 32'hf13629e9 ;
    mem[8'ha8] <= 32'hd0b3ba59 ;
    mem[8'ha9] <= 32'hd6ff9389 ;
    mem[8'haa] <= 32'hdc2be9f9 ;
    mem[8'hab] <= 32'hda67c029 ;
    mem[8'hac] <= 32'hc9831d19 ;
    mem[8'had] <= 32'hcfcf34c9 ;
    mem[8'hae] <= 32'hc51b4eb9 ;
    mem[8'haf] <= 32'hc3576769 ;
    mem[8'hb0] <= 32'h861069d9 ;
    mem[8'hb1] <= 32'h805c4009 ;
    mem[8'hb2] <= 32'h8a883a79 ;
    mem[8'hb3] <= 32'h8cc413a9 ;
    mem[8'hb4] <= 32'h9f20ce99 ;
    mem[8'hb5] <= 32'h996ce749 ;
    mem[8'hb6] <= 32'h93b89d39 ;
    mem[8'hb7] <= 32'h95f4b4e9 ;
    mem[8'hb8] <= 32'hb4712759 ;
    mem[8'hb9] <= 32'hb23d0e89 ;
    mem[8'hba] <= 32'hb8e974f9 ;
    mem[8'hbb] <= 32'hbea55d29 ;
    mem[8'hbc] <= 32'had418019 ;
    mem[8'hbd] <= 32'hab0da9c9 ;
    mem[8'hbe] <= 32'ha1d9d3b9 ;
    mem[8'hbf] <= 32'ha795fa69 ;
    mem[8'hc0] <= 32'hbc9ca76e ;
    mem[8'hc1] <= 32'hbad08ebe ;
    mem[8'hc2] <= 32'hb004f4ce ;
    mem[8'hc3] <= 32'hb648dd1e ;
    mem[8'hc4] <= 32'ha5ac002e ;
    mem[8'hc5] <= 32'ha3e029fe ;
    mem[8'hc6] <= 32'ha934538e ;
    mem[8'hc7] <= 32'haf787a5e ;
    mem[8'hc8] <= 32'h8efde9ee ;
    mem[8'hc9] <= 32'h88b1c03e ;
    mem[8'hca] <= 32'h8265ba4e ;
    mem[8'hcb] <= 32'h8429939e ;
    mem[8'hcc] <= 32'h97cd4eae ;
    mem[8'hcd] <= 32'h9181677e ;
    mem[8'hce] <= 32'h9b551d0e ;
    mem[8'hcf] <= 32'h9d1934de ;
    mem[8'hd0] <= 32'hd85e3a6e ;
    mem[8'hd1] <= 32'hde1213be ;
    mem[8'hd2] <= 32'hd4c669ce ;
    mem[8'hd3] <= 32'hd28a401e ;
    mem[8'hd4] <= 32'hc16e9d2e ;
    mem[8'hd5] <= 32'hc722b4fe ;
    mem[8'hd6] <= 32'hcdf6ce8e ;
    mem[8'hd7] <= 32'hcbbae75e ;
    mem[8'hd8] <= 32'hea3f74ee ;
    mem[8'hd9] <= 32'hec735d3e ;
    mem[8'hda] <= 32'he6a7274e ;
    mem[8'hdb] <= 32'he0eb0e9e ;
    mem[8'hdc] <= 32'hf30fd3ae ;
    mem[8'hdd] <= 32'hf543fa7e ;
    mem[8'hde] <= 32'hff97800e ;
    mem[8'hdf] <= 32'hf9dba9de ;
    mem[8'he0] <= 32'h75199d6e ;
    mem[8'he1] <= 32'h7355b4be ;
    mem[8'he2] <= 32'h7981cece ;
    mem[8'he3] <= 32'h7fcde71e ;
    mem[8'he4] <= 32'h6c293a2e ;
    mem[8'he5] <= 32'h6a6513fe ;
    mem[8'he6] <= 32'h60b1698e ;
    mem[8'he7] <= 32'h66fd405e ;
    mem[8'he8] <= 32'h4778d3ee ;
    mem[8'he9] <= 32'h4134fa3e ;
    mem[8'hea] <= 32'h4be0804e ;
    mem[8'heb] <= 32'h4daca99e ;
    mem[8'hec] <= 32'h5e4874ae ;
    mem[8'hed] <= 32'h58045d7e ;
    mem[8'hee] <= 32'h52d0270e ;
    mem[8'hef] <= 32'h549c0ede ;
    mem[8'hf0] <= 32'h11db006e ;
    mem[8'hf1] <= 32'h179729be ;
    mem[8'hf2] <= 32'h1d4353ce ;
    mem[8'hf3] <= 32'h1b0f7a1e ;
    mem[8'hf4] <= 32'h8eba72e ;
    mem[8'hf5] <= 32'hea78efe ;
    mem[8'hf6] <= 32'h473f48e ;
    mem[8'hf7] <= 32'h23fdd5e ;
    mem[8'hf8] <= 32'h23ba4eee ;
    mem[8'hf9] <= 32'h25f6673e ;
    mem[8'hfa] <= 32'h2f221d4e ;
    mem[8'hfb] <= 32'h296e349e ;
    mem[8'hfc] <= 32'h3a8ae9ae ;
    mem[8'hfd] <= 32'h3cc6c07e ;
    mem[8'hfe] <= 32'h3612ba0e ;
    mem[8'hff] <= 32'h305e93de ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
