module crctab_ev12
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'he8a45605 ;
    mem[8'h2] <= 32'hd589b1bd ;
    mem[8'h3] <= 32'h3d2de7b8 ;
    mem[8'h4] <= 32'hafd27ecd ;
    mem[8'h5] <= 32'h477628c8 ;
    mem[8'h6] <= 32'h7a5bcf70 ;
    mem[8'h7] <= 32'h92ff9975 ;
    mem[8'h8] <= 32'h5b65e02d ;
    mem[8'h9] <= 32'hb3c1b628 ;
    mem[8'ha] <= 32'h8eec5190 ;
    mem[8'hb] <= 32'h66480795 ;
    mem[8'hc] <= 32'hf4b79ee0 ;
    mem[8'hd] <= 32'h1c13c8e5 ;
    mem[8'he] <= 32'h213e2f5d ;
    mem[8'hf] <= 32'hc99a7958 ;
    mem[8'h10] <= 32'hb6cbc05a ;
    mem[8'h11] <= 32'h5e6f965f ;
    mem[8'h12] <= 32'h634271e7 ;
    mem[8'h13] <= 32'h8be627e2 ;
    mem[8'h14] <= 32'h1919be97 ;
    mem[8'h15] <= 32'hf1bde892 ;
    mem[8'h16] <= 32'hcc900f2a ;
    mem[8'h17] <= 32'h2434592f ;
    mem[8'h18] <= 32'hedae2077 ;
    mem[8'h19] <= 32'h50a7672 ;
    mem[8'h1a] <= 32'h382791ca ;
    mem[8'h1b] <= 32'hd083c7cf ;
    mem[8'h1c] <= 32'h427c5eba ;
    mem[8'h1d] <= 32'haad808bf ;
    mem[8'h1e] <= 32'h97f5ef07 ;
    mem[8'h1f] <= 32'h7f51b902 ;
    mem[8'h20] <= 32'h69569d03 ;
    mem[8'h21] <= 32'h81f2cb06 ;
    mem[8'h22] <= 32'hbcdf2cbe ;
    mem[8'h23] <= 32'h547b7abb ;
    mem[8'h24] <= 32'hc684e3ce ;
    mem[8'h25] <= 32'h2e20b5cb ;
    mem[8'h26] <= 32'h130d5273 ;
    mem[8'h27] <= 32'hfba90476 ;
    mem[8'h28] <= 32'h32337d2e ;
    mem[8'h29] <= 32'hda972b2b ;
    mem[8'h2a] <= 32'he7bacc93 ;
    mem[8'h2b] <= 32'hf1e9a96 ;
    mem[8'h2c] <= 32'h9de103e3 ;
    mem[8'h2d] <= 32'h754555e6 ;
    mem[8'h2e] <= 32'h4868b25e ;
    mem[8'h2f] <= 32'ha0cce45b ;
    mem[8'h30] <= 32'hdf9d5d59 ;
    mem[8'h31] <= 32'h37390b5c ;
    mem[8'h32] <= 32'ha14ece4 ;
    mem[8'h33] <= 32'he2b0bae1 ;
    mem[8'h34] <= 32'h704f2394 ;
    mem[8'h35] <= 32'h98eb7591 ;
    mem[8'h36] <= 32'ha5c69229 ;
    mem[8'h37] <= 32'h4d62c42c ;
    mem[8'h38] <= 32'h84f8bd74 ;
    mem[8'h39] <= 32'h6c5ceb71 ;
    mem[8'h3a] <= 32'h51710cc9 ;
    mem[8'h3b] <= 32'hb9d55acc ;
    mem[8'h3c] <= 32'h2b2ac3b9 ;
    mem[8'h3d] <= 32'hc38e95bc ;
    mem[8'h3e] <= 32'hfea37204 ;
    mem[8'h3f] <= 32'h16072401 ;
    mem[8'h40] <= 32'hd2ad3a06 ;
    mem[8'h41] <= 32'h3a096c03 ;
    mem[8'h42] <= 32'h7248bbb ;
    mem[8'h43] <= 32'hef80ddbe ;
    mem[8'h44] <= 32'h7d7f44cb ;
    mem[8'h45] <= 32'h95db12ce ;
    mem[8'h46] <= 32'ha8f6f576 ;
    mem[8'h47] <= 32'h4052a373 ;
    mem[8'h48] <= 32'h89c8da2b ;
    mem[8'h49] <= 32'h616c8c2e ;
    mem[8'h4a] <= 32'h5c416b96 ;
    mem[8'h4b] <= 32'hb4e53d93 ;
    mem[8'h4c] <= 32'h261aa4e6 ;
    mem[8'h4d] <= 32'hcebef2e3 ;
    mem[8'h4e] <= 32'hf393155b ;
    mem[8'h4f] <= 32'h1b37435e ;
    mem[8'h50] <= 32'h6466fa5c ;
    mem[8'h51] <= 32'h8cc2ac59 ;
    mem[8'h52] <= 32'hb1ef4be1 ;
    mem[8'h53] <= 32'h594b1de4 ;
    mem[8'h54] <= 32'hcbb48491 ;
    mem[8'h55] <= 32'h2310d294 ;
    mem[8'h56] <= 32'h1e3d352c ;
    mem[8'h57] <= 32'hf6996329 ;
    mem[8'h58] <= 32'h3f031a71 ;
    mem[8'h59] <= 32'hd7a74c74 ;
    mem[8'h5a] <= 32'hea8aabcc ;
    mem[8'h5b] <= 32'h22efdc9 ;
    mem[8'h5c] <= 32'h90d164bc ;
    mem[8'h5d] <= 32'h787532b9 ;
    mem[8'h5e] <= 32'h4558d501 ;
    mem[8'h5f] <= 32'hadfc8304 ;
    mem[8'h60] <= 32'hbbfba705 ;
    mem[8'h61] <= 32'h535ff100 ;
    mem[8'h62] <= 32'h6e7216b8 ;
    mem[8'h63] <= 32'h86d640bd ;
    mem[8'h64] <= 32'h1429d9c8 ;
    mem[8'h65] <= 32'hfc8d8fcd ;
    mem[8'h66] <= 32'hc1a06875 ;
    mem[8'h67] <= 32'h29043e70 ;
    mem[8'h68] <= 32'he09e4728 ;
    mem[8'h69] <= 32'h83a112d ;
    mem[8'h6a] <= 32'h3517f695 ;
    mem[8'h6b] <= 32'hddb3a090 ;
    mem[8'h6c] <= 32'h4f4c39e5 ;
    mem[8'h6d] <= 32'ha7e86fe0 ;
    mem[8'h6e] <= 32'h9ac58858 ;
    mem[8'h6f] <= 32'h7261de5d ;
    mem[8'h70] <= 32'hd30675f ;
    mem[8'h71] <= 32'he594315a ;
    mem[8'h72] <= 32'hd8b9d6e2 ;
    mem[8'h73] <= 32'h301d80e7 ;
    mem[8'h74] <= 32'ha2e21992 ;
    mem[8'h75] <= 32'h4a464f97 ;
    mem[8'h76] <= 32'h776ba82f ;
    mem[8'h77] <= 32'h9fcffe2a ;
    mem[8'h78] <= 32'h56558772 ;
    mem[8'h79] <= 32'hbef1d177 ;
    mem[8'h7a] <= 32'h83dc36cf ;
    mem[8'h7b] <= 32'h6b7860ca ;
    mem[8'h7c] <= 32'hf987f9bf ;
    mem[8'h7d] <= 32'h1123afba ;
    mem[8'h7e] <= 32'h2c0e4802 ;
    mem[8'h7f] <= 32'hc4aa1e07 ;
    mem[8'h80] <= 32'ha19b69bb ;
    mem[8'h81] <= 32'h493f3fbe ;
    mem[8'h82] <= 32'h7412d806 ;
    mem[8'h83] <= 32'h9cb68e03 ;
    mem[8'h84] <= 32'he491776 ;
    mem[8'h85] <= 32'he6ed4173 ;
    mem[8'h86] <= 32'hdbc0a6cb ;
    mem[8'h87] <= 32'h3364f0ce ;
    mem[8'h88] <= 32'hfafe8996 ;
    mem[8'h89] <= 32'h125adf93 ;
    mem[8'h8a] <= 32'h2f77382b ;
    mem[8'h8b] <= 32'hc7d36e2e ;
    mem[8'h8c] <= 32'h552cf75b ;
    mem[8'h8d] <= 32'hbd88a15e ;
    mem[8'h8e] <= 32'h80a546e6 ;
    mem[8'h8f] <= 32'h680110e3 ;
    mem[8'h90] <= 32'h1750a9e1 ;
    mem[8'h91] <= 32'hfff4ffe4 ;
    mem[8'h92] <= 32'hc2d9185c ;
    mem[8'h93] <= 32'h2a7d4e59 ;
    mem[8'h94] <= 32'hb882d72c ;
    mem[8'h95] <= 32'h50268129 ;
    mem[8'h96] <= 32'h6d0b6691 ;
    mem[8'h97] <= 32'h85af3094 ;
    mem[8'h98] <= 32'h4c3549cc ;
    mem[8'h99] <= 32'ha4911fc9 ;
    mem[8'h9a] <= 32'h99bcf871 ;
    mem[8'h9b] <= 32'h7118ae74 ;
    mem[8'h9c] <= 32'he3e73701 ;
    mem[8'h9d] <= 32'hb436104 ;
    mem[8'h9e] <= 32'h366e86bc ;
    mem[8'h9f] <= 32'hdecad0b9 ;
    mem[8'ha0] <= 32'hc8cdf4b8 ;
    mem[8'ha1] <= 32'h2069a2bd ;
    mem[8'ha2] <= 32'h1d444505 ;
    mem[8'ha3] <= 32'hf5e01300 ;
    mem[8'ha4] <= 32'h671f8a75 ;
    mem[8'ha5] <= 32'h8fbbdc70 ;
    mem[8'ha6] <= 32'hb2963bc8 ;
    mem[8'ha7] <= 32'h5a326dcd ;
    mem[8'ha8] <= 32'h93a81495 ;
    mem[8'ha9] <= 32'h7b0c4290 ;
    mem[8'haa] <= 32'h4621a528 ;
    mem[8'hab] <= 32'hae85f32d ;
    mem[8'hac] <= 32'h3c7a6a58 ;
    mem[8'had] <= 32'hd4de3c5d ;
    mem[8'hae] <= 32'he9f3dbe5 ;
    mem[8'haf] <= 32'h1578de0 ;
    mem[8'hb0] <= 32'h7e0634e2 ;
    mem[8'hb1] <= 32'h96a262e7 ;
    mem[8'hb2] <= 32'hab8f855f ;
    mem[8'hb3] <= 32'h432bd35a ;
    mem[8'hb4] <= 32'hd1d44a2f ;
    mem[8'hb5] <= 32'h39701c2a ;
    mem[8'hb6] <= 32'h45dfb92 ;
    mem[8'hb7] <= 32'hecf9ad97 ;
    mem[8'hb8] <= 32'h2563d4cf ;
    mem[8'hb9] <= 32'hcdc782ca ;
    mem[8'hba] <= 32'hf0ea6572 ;
    mem[8'hbb] <= 32'h184e3377 ;
    mem[8'hbc] <= 32'h8ab1aa02 ;
    mem[8'hbd] <= 32'h6215fc07 ;
    mem[8'hbe] <= 32'h5f381bbf ;
    mem[8'hbf] <= 32'hb79c4dba ;
    mem[8'hc0] <= 32'h733653bd ;
    mem[8'hc1] <= 32'h9b9205b8 ;
    mem[8'hc2] <= 32'ha6bfe200 ;
    mem[8'hc3] <= 32'h4e1bb405 ;
    mem[8'hc4] <= 32'hdce42d70 ;
    mem[8'hc5] <= 32'h34407b75 ;
    mem[8'hc6] <= 32'h96d9ccd ;
    mem[8'hc7] <= 32'he1c9cac8 ;
    mem[8'hc8] <= 32'h2853b390 ;
    mem[8'hc9] <= 32'hc0f7e595 ;
    mem[8'hca] <= 32'hfdda022d ;
    mem[8'hcb] <= 32'h157e5428 ;
    mem[8'hcc] <= 32'h8781cd5d ;
    mem[8'hcd] <= 32'h6f259b58 ;
    mem[8'hce] <= 32'h52087ce0 ;
    mem[8'hcf] <= 32'hbaac2ae5 ;
    mem[8'hd0] <= 32'hc5fd93e7 ;
    mem[8'hd1] <= 32'h2d59c5e2 ;
    mem[8'hd2] <= 32'h1074225a ;
    mem[8'hd3] <= 32'hf8d0745f ;
    mem[8'hd4] <= 32'h6a2fed2a ;
    mem[8'hd5] <= 32'h828bbb2f ;
    mem[8'hd6] <= 32'hbfa65c97 ;
    mem[8'hd7] <= 32'h57020a92 ;
    mem[8'hd8] <= 32'h9e9873ca ;
    mem[8'hd9] <= 32'h763c25cf ;
    mem[8'hda] <= 32'h4b11c277 ;
    mem[8'hdb] <= 32'ha3b59472 ;
    mem[8'hdc] <= 32'h314a0d07 ;
    mem[8'hdd] <= 32'hd9ee5b02 ;
    mem[8'hde] <= 32'he4c3bcba ;
    mem[8'hdf] <= 32'hc67eabf ;
    mem[8'he0] <= 32'h1a60cebe ;
    mem[8'he1] <= 32'hf2c498bb ;
    mem[8'he2] <= 32'hcfe97f03 ;
    mem[8'he3] <= 32'h274d2906 ;
    mem[8'he4] <= 32'hb5b2b073 ;
    mem[8'he5] <= 32'h5d16e676 ;
    mem[8'he6] <= 32'h603b01ce ;
    mem[8'he7] <= 32'h889f57cb ;
    mem[8'he8] <= 32'h41052e93 ;
    mem[8'he9] <= 32'ha9a17896 ;
    mem[8'hea] <= 32'h948c9f2e ;
    mem[8'heb] <= 32'h7c28c92b ;
    mem[8'hec] <= 32'heed7505e ;
    mem[8'hed] <= 32'h673065b ;
    mem[8'hee] <= 32'h3b5ee1e3 ;
    mem[8'hef] <= 32'hd3fab7e6 ;
    mem[8'hf0] <= 32'hacab0ee4 ;
    mem[8'hf1] <= 32'h440f58e1 ;
    mem[8'hf2] <= 32'h7922bf59 ;
    mem[8'hf3] <= 32'h9186e95c ;
    mem[8'hf4] <= 32'h3797029 ;
    mem[8'hf5] <= 32'hebdd262c ;
    mem[8'hf6] <= 32'hd6f0c194 ;
    mem[8'hf7] <= 32'h3e549791 ;
    mem[8'hf8] <= 32'hf7ceeec9 ;
    mem[8'hf9] <= 32'h1f6ab8cc ;
    mem[8'hfa] <= 32'h22475f74 ;
    mem[8'hfb] <= 32'hcae30971 ;
    mem[8'hfc] <= 32'h581c9004 ;
    mem[8'hfd] <= 32'hb0b8c601 ;
    mem[8'hfe] <= 32'h8d9521b9 ;
    mem[8'hff] <= 32'h653177bc ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
