module crctab_ev5
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h1b280d78 ;
    mem[8'h2] <= 32'h36501af0 ;
    mem[8'h3] <= 32'h2d781788 ;
    mem[8'h4] <= 32'h6ca035e0 ;
    mem[8'h5] <= 32'h77883898 ;
    mem[8'h6] <= 32'h5af02f10 ;
    mem[8'h7] <= 32'h41d82268 ;
    mem[8'h8] <= 32'hd9406bc0 ;
    mem[8'h9] <= 32'hc26866b8 ;
    mem[8'ha] <= 32'hef107130 ;
    mem[8'hb] <= 32'hf4387c48 ;
    mem[8'hc] <= 32'hb5e05e20 ;
    mem[8'hd] <= 32'haec85358 ;
    mem[8'he] <= 32'h83b044d0 ;
    mem[8'hf] <= 32'h989849a8 ;
    mem[8'h10] <= 32'hb641ca37 ;
    mem[8'h11] <= 32'had69c74f ;
    mem[8'h12] <= 32'h8011d0c7 ;
    mem[8'h13] <= 32'h9b39ddbf ;
    mem[8'h14] <= 32'hdae1ffd7 ;
    mem[8'h15] <= 32'hc1c9f2af ;
    mem[8'h16] <= 32'hecb1e527 ;
    mem[8'h17] <= 32'hf799e85f ;
    mem[8'h18] <= 32'h6f01a1f7 ;
    mem[8'h19] <= 32'h7429ac8f ;
    mem[8'h1a] <= 32'h5951bb07 ;
    mem[8'h1b] <= 32'h4279b67f ;
    mem[8'h1c] <= 32'h3a19417 ;
    mem[8'h1d] <= 32'h1889996f ;
    mem[8'h1e] <= 32'h35f18ee7 ;
    mem[8'h1f] <= 32'h2ed9839f ;
    mem[8'h20] <= 32'h684289d9 ;
    mem[8'h21] <= 32'h736a84a1 ;
    mem[8'h22] <= 32'h5e129329 ;
    mem[8'h23] <= 32'h453a9e51 ;
    mem[8'h24] <= 32'h4e2bc39 ;
    mem[8'h25] <= 32'h1fcab141 ;
    mem[8'h26] <= 32'h32b2a6c9 ;
    mem[8'h27] <= 32'h299aabb1 ;
    mem[8'h28] <= 32'hb102e219 ;
    mem[8'h29] <= 32'haa2aef61 ;
    mem[8'h2a] <= 32'h8752f8e9 ;
    mem[8'h2b] <= 32'h9c7af591 ;
    mem[8'h2c] <= 32'hdda2d7f9 ;
    mem[8'h2d] <= 32'hc68ada81 ;
    mem[8'h2e] <= 32'hebf2cd09 ;
    mem[8'h2f] <= 32'hf0dac071 ;
    mem[8'h30] <= 32'hde0343ee ;
    mem[8'h31] <= 32'hc52b4e96 ;
    mem[8'h32] <= 32'he853591e ;
    mem[8'h33] <= 32'hf37b5466 ;
    mem[8'h34] <= 32'hb2a3760e ;
    mem[8'h35] <= 32'ha98b7b76 ;
    mem[8'h36] <= 32'h84f36cfe ;
    mem[8'h37] <= 32'h9fdb6186 ;
    mem[8'h38] <= 32'h743282e ;
    mem[8'h39] <= 32'h1c6b2556 ;
    mem[8'h3a] <= 32'h311332de ;
    mem[8'h3b] <= 32'h2a3b3fa6 ;
    mem[8'h3c] <= 32'h6be31dce ;
    mem[8'h3d] <= 32'h70cb10b6 ;
    mem[8'h3e] <= 32'h5db3073e ;
    mem[8'h3f] <= 32'h469b0a46 ;
    mem[8'h40] <= 32'hd08513b2 ;
    mem[8'h41] <= 32'hcbad1eca ;
    mem[8'h42] <= 32'he6d50942 ;
    mem[8'h43] <= 32'hfdfd043a ;
    mem[8'h44] <= 32'hbc252652 ;
    mem[8'h45] <= 32'ha70d2b2a ;
    mem[8'h46] <= 32'h8a753ca2 ;
    mem[8'h47] <= 32'h915d31da ;
    mem[8'h48] <= 32'h9c57872 ;
    mem[8'h49] <= 32'h12ed750a ;
    mem[8'h4a] <= 32'h3f956282 ;
    mem[8'h4b] <= 32'h24bd6ffa ;
    mem[8'h4c] <= 32'h65654d92 ;
    mem[8'h4d] <= 32'h7e4d40ea ;
    mem[8'h4e] <= 32'h53355762 ;
    mem[8'h4f] <= 32'h481d5a1a ;
    mem[8'h50] <= 32'h66c4d985 ;
    mem[8'h51] <= 32'h7decd4fd ;
    mem[8'h52] <= 32'h5094c375 ;
    mem[8'h53] <= 32'h4bbcce0d ;
    mem[8'h54] <= 32'ha64ec65 ;
    mem[8'h55] <= 32'h114ce11d ;
    mem[8'h56] <= 32'h3c34f695 ;
    mem[8'h57] <= 32'h271cfbed ;
    mem[8'h58] <= 32'hbf84b245 ;
    mem[8'h59] <= 32'ha4acbf3d ;
    mem[8'h5a] <= 32'h89d4a8b5 ;
    mem[8'h5b] <= 32'h92fca5cd ;
    mem[8'h5c] <= 32'hd32487a5 ;
    mem[8'h5d] <= 32'hc80c8add ;
    mem[8'h5e] <= 32'he5749d55 ;
    mem[8'h5f] <= 32'hfe5c902d ;
    mem[8'h60] <= 32'hb8c79a6b ;
    mem[8'h61] <= 32'ha3ef9713 ;
    mem[8'h62] <= 32'h8e97809b ;
    mem[8'h63] <= 32'h95bf8de3 ;
    mem[8'h64] <= 32'hd467af8b ;
    mem[8'h65] <= 32'hcf4fa2f3 ;
    mem[8'h66] <= 32'he237b57b ;
    mem[8'h67] <= 32'hf91fb803 ;
    mem[8'h68] <= 32'h6187f1ab ;
    mem[8'h69] <= 32'h7aaffcd3 ;
    mem[8'h6a] <= 32'h57d7eb5b ;
    mem[8'h6b] <= 32'h4cffe623 ;
    mem[8'h6c] <= 32'hd27c44b ;
    mem[8'h6d] <= 32'h160fc933 ;
    mem[8'h6e] <= 32'h3b77debb ;
    mem[8'h6f] <= 32'h205fd3c3 ;
    mem[8'h70] <= 32'he86505c ;
    mem[8'h71] <= 32'h15ae5d24 ;
    mem[8'h72] <= 32'h38d64aac ;
    mem[8'h73] <= 32'h23fe47d4 ;
    mem[8'h74] <= 32'h622665bc ;
    mem[8'h75] <= 32'h790e68c4 ;
    mem[8'h76] <= 32'h54767f4c ;
    mem[8'h77] <= 32'h4f5e7234 ;
    mem[8'h78] <= 32'hd7c63b9c ;
    mem[8'h79] <= 32'hccee36e4 ;
    mem[8'h7a] <= 32'he196216c ;
    mem[8'h7b] <= 32'hfabe2c14 ;
    mem[8'h7c] <= 32'hbb660e7c ;
    mem[8'h7d] <= 32'ha04e0304 ;
    mem[8'h7e] <= 32'h8d36148c ;
    mem[8'h7f] <= 32'h961e19f4 ;
    mem[8'h80] <= 32'ha5cb3ad3 ;
    mem[8'h81] <= 32'hbee337ab ;
    mem[8'h82] <= 32'h939b2023 ;
    mem[8'h83] <= 32'h88b32d5b ;
    mem[8'h84] <= 32'hc96b0f33 ;
    mem[8'h85] <= 32'hd243024b ;
    mem[8'h86] <= 32'hff3b15c3 ;
    mem[8'h87] <= 32'he41318bb ;
    mem[8'h88] <= 32'h7c8b5113 ;
    mem[8'h89] <= 32'h67a35c6b ;
    mem[8'h8a] <= 32'h4adb4be3 ;
    mem[8'h8b] <= 32'h51f3469b ;
    mem[8'h8c] <= 32'h102b64f3 ;
    mem[8'h8d] <= 32'hb03698b ;
    mem[8'h8e] <= 32'h267b7e03 ;
    mem[8'h8f] <= 32'h3d53737b ;
    mem[8'h90] <= 32'h138af0e4 ;
    mem[8'h91] <= 32'h8a2fd9c ;
    mem[8'h92] <= 32'h25daea14 ;
    mem[8'h93] <= 32'h3ef2e76c ;
    mem[8'h94] <= 32'h7f2ac504 ;
    mem[8'h95] <= 32'h6402c87c ;
    mem[8'h96] <= 32'h497adff4 ;
    mem[8'h97] <= 32'h5252d28c ;
    mem[8'h98] <= 32'hcaca9b24 ;
    mem[8'h99] <= 32'hd1e2965c ;
    mem[8'h9a] <= 32'hfc9a81d4 ;
    mem[8'h9b] <= 32'he7b28cac ;
    mem[8'h9c] <= 32'ha66aaec4 ;
    mem[8'h9d] <= 32'hbd42a3bc ;
    mem[8'h9e] <= 32'h903ab434 ;
    mem[8'h9f] <= 32'h8b12b94c ;
    mem[8'ha0] <= 32'hcd89b30a ;
    mem[8'ha1] <= 32'hd6a1be72 ;
    mem[8'ha2] <= 32'hfbd9a9fa ;
    mem[8'ha3] <= 32'he0f1a482 ;
    mem[8'ha4] <= 32'ha12986ea ;
    mem[8'ha5] <= 32'hba018b92 ;
    mem[8'ha6] <= 32'h97799c1a ;
    mem[8'ha7] <= 32'h8c519162 ;
    mem[8'ha8] <= 32'h14c9d8ca ;
    mem[8'ha9] <= 32'hfe1d5b2 ;
    mem[8'haa] <= 32'h2299c23a ;
    mem[8'hab] <= 32'h39b1cf42 ;
    mem[8'hac] <= 32'h7869ed2a ;
    mem[8'had] <= 32'h6341e052 ;
    mem[8'hae] <= 32'h4e39f7da ;
    mem[8'haf] <= 32'h5511faa2 ;
    mem[8'hb0] <= 32'h7bc8793d ;
    mem[8'hb1] <= 32'h60e07445 ;
    mem[8'hb2] <= 32'h4d9863cd ;
    mem[8'hb3] <= 32'h56b06eb5 ;
    mem[8'hb4] <= 32'h17684cdd ;
    mem[8'hb5] <= 32'hc4041a5 ;
    mem[8'hb6] <= 32'h2138562d ;
    mem[8'hb7] <= 32'h3a105b55 ;
    mem[8'hb8] <= 32'ha28812fd ;
    mem[8'hb9] <= 32'hb9a01f85 ;
    mem[8'hba] <= 32'h94d8080d ;
    mem[8'hbb] <= 32'h8ff00575 ;
    mem[8'hbc] <= 32'hce28271d ;
    mem[8'hbd] <= 32'hd5002a65 ;
    mem[8'hbe] <= 32'hf8783ded ;
    mem[8'hbf] <= 32'he3503095 ;
    mem[8'hc0] <= 32'h754e2961 ;
    mem[8'hc1] <= 32'h6e662419 ;
    mem[8'hc2] <= 32'h431e3391 ;
    mem[8'hc3] <= 32'h58363ee9 ;
    mem[8'hc4] <= 32'h19ee1c81 ;
    mem[8'hc5] <= 32'h2c611f9 ;
    mem[8'hc6] <= 32'h2fbe0671 ;
    mem[8'hc7] <= 32'h34960b09 ;
    mem[8'hc8] <= 32'hac0e42a1 ;
    mem[8'hc9] <= 32'hb7264fd9 ;
    mem[8'hca] <= 32'h9a5e5851 ;
    mem[8'hcb] <= 32'h81765529 ;
    mem[8'hcc] <= 32'hc0ae7741 ;
    mem[8'hcd] <= 32'hdb867a39 ;
    mem[8'hce] <= 32'hf6fe6db1 ;
    mem[8'hcf] <= 32'hedd660c9 ;
    mem[8'hd0] <= 32'hc30fe356 ;
    mem[8'hd1] <= 32'hd827ee2e ;
    mem[8'hd2] <= 32'hf55ff9a6 ;
    mem[8'hd3] <= 32'hee77f4de ;
    mem[8'hd4] <= 32'hafafd6b6 ;
    mem[8'hd5] <= 32'hb487dbce ;
    mem[8'hd6] <= 32'h99ffcc46 ;
    mem[8'hd7] <= 32'h82d7c13e ;
    mem[8'hd8] <= 32'h1a4f8896 ;
    mem[8'hd9] <= 32'h16785ee ;
    mem[8'hda] <= 32'h2c1f9266 ;
    mem[8'hdb] <= 32'h37379f1e ;
    mem[8'hdc] <= 32'h76efbd76 ;
    mem[8'hdd] <= 32'h6dc7b00e ;
    mem[8'hde] <= 32'h40bfa786 ;
    mem[8'hdf] <= 32'h5b97aafe ;
    mem[8'he0] <= 32'h1d0ca0b8 ;
    mem[8'he1] <= 32'h624adc0 ;
    mem[8'he2] <= 32'h2b5cba48 ;
    mem[8'he3] <= 32'h3074b730 ;
    mem[8'he4] <= 32'h71ac9558 ;
    mem[8'he5] <= 32'h6a849820 ;
    mem[8'he6] <= 32'h47fc8fa8 ;
    mem[8'he7] <= 32'h5cd482d0 ;
    mem[8'he8] <= 32'hc44ccb78 ;
    mem[8'he9] <= 32'hdf64c600 ;
    mem[8'hea] <= 32'hf21cd188 ;
    mem[8'heb] <= 32'he934dcf0 ;
    mem[8'hec] <= 32'ha8ecfe98 ;
    mem[8'hed] <= 32'hb3c4f3e0 ;
    mem[8'hee] <= 32'h9ebce468 ;
    mem[8'hef] <= 32'h8594e910 ;
    mem[8'hf0] <= 32'hab4d6a8f ;
    mem[8'hf1] <= 32'hb06567f7 ;
    mem[8'hf2] <= 32'h9d1d707f ;
    mem[8'hf3] <= 32'h86357d07 ;
    mem[8'hf4] <= 32'hc7ed5f6f ;
    mem[8'hf5] <= 32'hdcc55217 ;
    mem[8'hf6] <= 32'hf1bd459f ;
    mem[8'hf7] <= 32'hea9548e7 ;
    mem[8'hf8] <= 32'h720d014f ;
    mem[8'hf9] <= 32'h69250c37 ;
    mem[8'hfa] <= 32'h445d1bbf ;
    mem[8'hfb] <= 32'h5f7516c7 ;
    mem[8'hfc] <= 32'h1ead34af ;
    mem[8'hfd] <= 32'h58539d7 ;
    mem[8'hfe] <= 32'h28fd2e5f ;
    mem[8'hff] <= 32'h33d52327 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
