module crctab_ev0
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h4c11db7 ;
    mem[8'h2] <= 32'h9823b6e ;
    mem[8'h3] <= 32'hd4326d9 ;
    mem[8'h4] <= 32'h130476dc ;
    mem[8'h5] <= 32'h17c56b6b ;
    mem[8'h6] <= 32'h1a864db2 ;
    mem[8'h7] <= 32'h1e475005 ;
    mem[8'h8] <= 32'h2608edb8 ;
    mem[8'h9] <= 32'h22c9f00f ;
    mem[8'ha] <= 32'h2f8ad6d6 ;
    mem[8'hb] <= 32'h2b4bcb61 ;
    mem[8'hc] <= 32'h350c9b64 ;
    mem[8'hd] <= 32'h31cd86d3 ;
    mem[8'he] <= 32'h3c8ea00a ;
    mem[8'hf] <= 32'h384fbdbd ;
    mem[8'h10] <= 32'h4c11db70 ;
    mem[8'h11] <= 32'h48d0c6c7 ;
    mem[8'h12] <= 32'h4593e01e ;
    mem[8'h13] <= 32'h4152fda9 ;
    mem[8'h14] <= 32'h5f15adac ;
    mem[8'h15] <= 32'h5bd4b01b ;
    mem[8'h16] <= 32'h569796c2 ;
    mem[8'h17] <= 32'h52568b75 ;
    mem[8'h18] <= 32'h6a1936c8 ;
    mem[8'h19] <= 32'h6ed82b7f ;
    mem[8'h1a] <= 32'h639b0da6 ;
    mem[8'h1b] <= 32'h675a1011 ;
    mem[8'h1c] <= 32'h791d4014 ;
    mem[8'h1d] <= 32'h7ddc5da3 ;
    mem[8'h1e] <= 32'h709f7b7a ;
    mem[8'h1f] <= 32'h745e66cd ;
    mem[8'h20] <= 32'h9823b6e0 ;
    mem[8'h21] <= 32'h9ce2ab57 ;
    mem[8'h22] <= 32'h91a18d8e ;
    mem[8'h23] <= 32'h95609039 ;
    mem[8'h24] <= 32'h8b27c03c ;
    mem[8'h25] <= 32'h8fe6dd8b ;
    mem[8'h26] <= 32'h82a5fb52 ;
    mem[8'h27] <= 32'h8664e6e5 ;
    mem[8'h28] <= 32'hbe2b5b58 ;
    mem[8'h29] <= 32'hbaea46ef ;
    mem[8'h2a] <= 32'hb7a96036 ;
    mem[8'h2b] <= 32'hb3687d81 ;
    mem[8'h2c] <= 32'had2f2d84 ;
    mem[8'h2d] <= 32'ha9ee3033 ;
    mem[8'h2e] <= 32'ha4ad16ea ;
    mem[8'h2f] <= 32'ha06c0b5d ;
    mem[8'h30] <= 32'hd4326d90 ;
    mem[8'h31] <= 32'hd0f37027 ;
    mem[8'h32] <= 32'hddb056fe ;
    mem[8'h33] <= 32'hd9714b49 ;
    mem[8'h34] <= 32'hc7361b4c ;
    mem[8'h35] <= 32'hc3f706fb ;
    mem[8'h36] <= 32'hceb42022 ;
    mem[8'h37] <= 32'hca753d95 ;
    mem[8'h38] <= 32'hf23a8028 ;
    mem[8'h39] <= 32'hf6fb9d9f ;
    mem[8'h3a] <= 32'hfbb8bb46 ;
    mem[8'h3b] <= 32'hff79a6f1 ;
    mem[8'h3c] <= 32'he13ef6f4 ;
    mem[8'h3d] <= 32'he5ffeb43 ;
    mem[8'h3e] <= 32'he8bccd9a ;
    mem[8'h3f] <= 32'hec7dd02d ;
    mem[8'h40] <= 32'h34867077 ;
    mem[8'h41] <= 32'h30476dc0 ;
    mem[8'h42] <= 32'h3d044b19 ;
    mem[8'h43] <= 32'h39c556ae ;
    mem[8'h44] <= 32'h278206ab ;
    mem[8'h45] <= 32'h23431b1c ;
    mem[8'h46] <= 32'h2e003dc5 ;
    mem[8'h47] <= 32'h2ac12072 ;
    mem[8'h48] <= 32'h128e9dcf ;
    mem[8'h49] <= 32'h164f8078 ;
    mem[8'h4a] <= 32'h1b0ca6a1 ;
    mem[8'h4b] <= 32'h1fcdbb16 ;
    mem[8'h4c] <= 32'h18aeb13 ;
    mem[8'h4d] <= 32'h54bf6a4 ;
    mem[8'h4e] <= 32'h808d07d ;
    mem[8'h4f] <= 32'hcc9cdca ;
    mem[8'h50] <= 32'h7897ab07 ;
    mem[8'h51] <= 32'h7c56b6b0 ;
    mem[8'h52] <= 32'h71159069 ;
    mem[8'h53] <= 32'h75d48dde ;
    mem[8'h54] <= 32'h6b93dddb ;
    mem[8'h55] <= 32'h6f52c06c ;
    mem[8'h56] <= 32'h6211e6b5 ;
    mem[8'h57] <= 32'h66d0fb02 ;
    mem[8'h58] <= 32'h5e9f46bf ;
    mem[8'h59] <= 32'h5a5e5b08 ;
    mem[8'h5a] <= 32'h571d7dd1 ;
    mem[8'h5b] <= 32'h53dc6066 ;
    mem[8'h5c] <= 32'h4d9b3063 ;
    mem[8'h5d] <= 32'h495a2dd4 ;
    mem[8'h5e] <= 32'h44190b0d ;
    mem[8'h5f] <= 32'h40d816ba ;
    mem[8'h60] <= 32'haca5c697 ;
    mem[8'h61] <= 32'ha864db20 ;
    mem[8'h62] <= 32'ha527fdf9 ;
    mem[8'h63] <= 32'ha1e6e04e ;
    mem[8'h64] <= 32'hbfa1b04b ;
    mem[8'h65] <= 32'hbb60adfc ;
    mem[8'h66] <= 32'hb6238b25 ;
    mem[8'h67] <= 32'hb2e29692 ;
    mem[8'h68] <= 32'h8aad2b2f ;
    mem[8'h69] <= 32'h8e6c3698 ;
    mem[8'h6a] <= 32'h832f1041 ;
    mem[8'h6b] <= 32'h87ee0df6 ;
    mem[8'h6c] <= 32'h99a95df3 ;
    mem[8'h6d] <= 32'h9d684044 ;
    mem[8'h6e] <= 32'h902b669d ;
    mem[8'h6f] <= 32'h94ea7b2a ;
    mem[8'h70] <= 32'he0b41de7 ;
    mem[8'h71] <= 32'he4750050 ;
    mem[8'h72] <= 32'he9362689 ;
    mem[8'h73] <= 32'hedf73b3e ;
    mem[8'h74] <= 32'hf3b06b3b ;
    mem[8'h75] <= 32'hf771768c ;
    mem[8'h76] <= 32'hfa325055 ;
    mem[8'h77] <= 32'hfef34de2 ;
    mem[8'h78] <= 32'hc6bcf05f ;
    mem[8'h79] <= 32'hc27dede8 ;
    mem[8'h7a] <= 32'hcf3ecb31 ;
    mem[8'h7b] <= 32'hcbffd686 ;
    mem[8'h7c] <= 32'hd5b88683 ;
    mem[8'h7d] <= 32'hd1799b34 ;
    mem[8'h7e] <= 32'hdc3abded ;
    mem[8'h7f] <= 32'hd8fba05a ;
    mem[8'h80] <= 32'h690ce0ee ;
    mem[8'h81] <= 32'h6dcdfd59 ;
    mem[8'h82] <= 32'h608edb80 ;
    mem[8'h83] <= 32'h644fc637 ;
    mem[8'h84] <= 32'h7a089632 ;
    mem[8'h85] <= 32'h7ec98b85 ;
    mem[8'h86] <= 32'h738aad5c ;
    mem[8'h87] <= 32'h774bb0eb ;
    mem[8'h88] <= 32'h4f040d56 ;
    mem[8'h89] <= 32'h4bc510e1 ;
    mem[8'h8a] <= 32'h46863638 ;
    mem[8'h8b] <= 32'h42472b8f ;
    mem[8'h8c] <= 32'h5c007b8a ;
    mem[8'h8d] <= 32'h58c1663d ;
    mem[8'h8e] <= 32'h558240e4 ;
    mem[8'h8f] <= 32'h51435d53 ;
    mem[8'h90] <= 32'h251d3b9e ;
    mem[8'h91] <= 32'h21dc2629 ;
    mem[8'h92] <= 32'h2c9f00f0 ;
    mem[8'h93] <= 32'h285e1d47 ;
    mem[8'h94] <= 32'h36194d42 ;
    mem[8'h95] <= 32'h32d850f5 ;
    mem[8'h96] <= 32'h3f9b762c ;
    mem[8'h97] <= 32'h3b5a6b9b ;
    mem[8'h98] <= 32'h315d626 ;
    mem[8'h99] <= 32'h7d4cb91 ;
    mem[8'h9a] <= 32'ha97ed48 ;
    mem[8'h9b] <= 32'he56f0ff ;
    mem[8'h9c] <= 32'h1011a0fa ;
    mem[8'h9d] <= 32'h14d0bd4d ;
    mem[8'h9e] <= 32'h19939b94 ;
    mem[8'h9f] <= 32'h1d528623 ;
    mem[8'ha0] <= 32'hf12f560e ;
    mem[8'ha1] <= 32'hf5ee4bb9 ;
    mem[8'ha2] <= 32'hf8ad6d60 ;
    mem[8'ha3] <= 32'hfc6c70d7 ;
    mem[8'ha4] <= 32'he22b20d2 ;
    mem[8'ha5] <= 32'he6ea3d65 ;
    mem[8'ha6] <= 32'heba91bbc ;
    mem[8'ha7] <= 32'hef68060b ;
    mem[8'ha8] <= 32'hd727bbb6 ;
    mem[8'ha9] <= 32'hd3e6a601 ;
    mem[8'haa] <= 32'hdea580d8 ;
    mem[8'hab] <= 32'hda649d6f ;
    mem[8'hac] <= 32'hc423cd6a ;
    mem[8'had] <= 32'hc0e2d0dd ;
    mem[8'hae] <= 32'hcda1f604 ;
    mem[8'haf] <= 32'hc960ebb3 ;
    mem[8'hb0] <= 32'hbd3e8d7e ;
    mem[8'hb1] <= 32'hb9ff90c9 ;
    mem[8'hb2] <= 32'hb4bcb610 ;
    mem[8'hb3] <= 32'hb07daba7 ;
    mem[8'hb4] <= 32'hae3afba2 ;
    mem[8'hb5] <= 32'haafbe615 ;
    mem[8'hb6] <= 32'ha7b8c0cc ;
    mem[8'hb7] <= 32'ha379dd7b ;
    mem[8'hb8] <= 32'h9b3660c6 ;
    mem[8'hb9] <= 32'h9ff77d71 ;
    mem[8'hba] <= 32'h92b45ba8 ;
    mem[8'hbb] <= 32'h9675461f ;
    mem[8'hbc] <= 32'h8832161a ;
    mem[8'hbd] <= 32'h8cf30bad ;
    mem[8'hbe] <= 32'h81b02d74 ;
    mem[8'hbf] <= 32'h857130c3 ;
    mem[8'hc0] <= 32'h5d8a9099 ;
    mem[8'hc1] <= 32'h594b8d2e ;
    mem[8'hc2] <= 32'h5408abf7 ;
    mem[8'hc3] <= 32'h50c9b640 ;
    mem[8'hc4] <= 32'h4e8ee645 ;
    mem[8'hc5] <= 32'h4a4ffbf2 ;
    mem[8'hc6] <= 32'h470cdd2b ;
    mem[8'hc7] <= 32'h43cdc09c ;
    mem[8'hc8] <= 32'h7b827d21 ;
    mem[8'hc9] <= 32'h7f436096 ;
    mem[8'hca] <= 32'h7200464f ;
    mem[8'hcb] <= 32'h76c15bf8 ;
    mem[8'hcc] <= 32'h68860bfd ;
    mem[8'hcd] <= 32'h6c47164a ;
    mem[8'hce] <= 32'h61043093 ;
    mem[8'hcf] <= 32'h65c52d24 ;
    mem[8'hd0] <= 32'h119b4be9 ;
    mem[8'hd1] <= 32'h155a565e ;
    mem[8'hd2] <= 32'h18197087 ;
    mem[8'hd3] <= 32'h1cd86d30 ;
    mem[8'hd4] <= 32'h29f3d35 ;
    mem[8'hd5] <= 32'h65e2082 ;
    mem[8'hd6] <= 32'hb1d065b ;
    mem[8'hd7] <= 32'hfdc1bec ;
    mem[8'hd8] <= 32'h3793a651 ;
    mem[8'hd9] <= 32'h3352bbe6 ;
    mem[8'hda] <= 32'h3e119d3f ;
    mem[8'hdb] <= 32'h3ad08088 ;
    mem[8'hdc] <= 32'h2497d08d ;
    mem[8'hdd] <= 32'h2056cd3a ;
    mem[8'hde] <= 32'h2d15ebe3 ;
    mem[8'hdf] <= 32'h29d4f654 ;
    mem[8'he0] <= 32'hc5a92679 ;
    mem[8'he1] <= 32'hc1683bce ;
    mem[8'he2] <= 32'hcc2b1d17 ;
    mem[8'he3] <= 32'hc8ea00a0 ;
    mem[8'he4] <= 32'hd6ad50a5 ;
    mem[8'he5] <= 32'hd26c4d12 ;
    mem[8'he6] <= 32'hdf2f6bcb ;
    mem[8'he7] <= 32'hdbee767c ;
    mem[8'he8] <= 32'he3a1cbc1 ;
    mem[8'he9] <= 32'he760d676 ;
    mem[8'hea] <= 32'hea23f0af ;
    mem[8'heb] <= 32'heee2ed18 ;
    mem[8'hec] <= 32'hf0a5bd1d ;
    mem[8'hed] <= 32'hf464a0aa ;
    mem[8'hee] <= 32'hf9278673 ;
    mem[8'hef] <= 32'hfde69bc4 ;
    mem[8'hf0] <= 32'h89b8fd09 ;
    mem[8'hf1] <= 32'h8d79e0be ;
    mem[8'hf2] <= 32'h803ac667 ;
    mem[8'hf3] <= 32'h84fbdbd0 ;
    mem[8'hf4] <= 32'h9abc8bd5 ;
    mem[8'hf5] <= 32'h9e7d9662 ;
    mem[8'hf6] <= 32'h933eb0bb ;
    mem[8'hf7] <= 32'h97ffad0c ;
    mem[8'hf8] <= 32'hafb010b1 ;
    mem[8'hf9] <= 32'hab710d06 ;
    mem[8'hfa] <= 32'ha6322bdf ;
    mem[8'hfb] <= 32'ha2f33668 ;
    mem[8'hfc] <= 32'hbcb4666d ;
    mem[8'hfd] <= 32'hb8757bda ;
    mem[8'hfe] <= 32'hb5365d03 ;
    mem[8'hff] <= 32'hb1f740b4 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
