module crctab_ev6
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h4f576811 ;
    mem[8'h2] <= 32'h9eaed022 ;
    mem[8'h3] <= 32'hd1f9b833 ;
    mem[8'h4] <= 32'h399cbdf3 ;
    mem[8'h5] <= 32'h76cbd5e2 ;
    mem[8'h6] <= 32'ha7326dd1 ;
    mem[8'h7] <= 32'he86505c0 ;
    mem[8'h8] <= 32'h73397be6 ;
    mem[8'h9] <= 32'h3c6e13f7 ;
    mem[8'ha] <= 32'hed97abc4 ;
    mem[8'hb] <= 32'ha2c0c3d5 ;
    mem[8'hc] <= 32'h4aa5c615 ;
    mem[8'hd] <= 32'h5f2ae04 ;
    mem[8'he] <= 32'hd40b1637 ;
    mem[8'hf] <= 32'h9b5c7e26 ;
    mem[8'h10] <= 32'he672f7cc ;
    mem[8'h11] <= 32'ha9259fdd ;
    mem[8'h12] <= 32'h78dc27ee ;
    mem[8'h13] <= 32'h378b4fff ;
    mem[8'h14] <= 32'hdfee4a3f ;
    mem[8'h15] <= 32'h90b9222e ;
    mem[8'h16] <= 32'h41409a1d ;
    mem[8'h17] <= 32'he17f20c ;
    mem[8'h18] <= 32'h954b8c2a ;
    mem[8'h19] <= 32'hda1ce43b ;
    mem[8'h1a] <= 32'hbe55c08 ;
    mem[8'h1b] <= 32'h44b23419 ;
    mem[8'h1c] <= 32'hacd731d9 ;
    mem[8'h1d] <= 32'he38059c8 ;
    mem[8'h1e] <= 32'h3279e1fb ;
    mem[8'h1f] <= 32'h7d2e89ea ;
    mem[8'h20] <= 32'hc824f22f ;
    mem[8'h21] <= 32'h87739a3e ;
    mem[8'h22] <= 32'h568a220d ;
    mem[8'h23] <= 32'h19dd4a1c ;
    mem[8'h24] <= 32'hf1b84fdc ;
    mem[8'h25] <= 32'hbeef27cd ;
    mem[8'h26] <= 32'h6f169ffe ;
    mem[8'h27] <= 32'h2041f7ef ;
    mem[8'h28] <= 32'hbb1d89c9 ;
    mem[8'h29] <= 32'hf44ae1d8 ;
    mem[8'h2a] <= 32'h25b359eb ;
    mem[8'h2b] <= 32'h6ae431fa ;
    mem[8'h2c] <= 32'h8281343a ;
    mem[8'h2d] <= 32'hcdd65c2b ;
    mem[8'h2e] <= 32'h1c2fe418 ;
    mem[8'h2f] <= 32'h53788c09 ;
    mem[8'h30] <= 32'h2e5605e3 ;
    mem[8'h31] <= 32'h61016df2 ;
    mem[8'h32] <= 32'hb0f8d5c1 ;
    mem[8'h33] <= 32'hffafbdd0 ;
    mem[8'h34] <= 32'h17cab810 ;
    mem[8'h35] <= 32'h589dd001 ;
    mem[8'h36] <= 32'h89646832 ;
    mem[8'h37] <= 32'hc6330023 ;
    mem[8'h38] <= 32'h5d6f7e05 ;
    mem[8'h39] <= 32'h12381614 ;
    mem[8'h3a] <= 32'hc3c1ae27 ;
    mem[8'h3b] <= 32'h8c96c636 ;
    mem[8'h3c] <= 32'h64f3c3f6 ;
    mem[8'h3d] <= 32'h2ba4abe7 ;
    mem[8'h3e] <= 32'hfa5d13d4 ;
    mem[8'h3f] <= 32'hb50a7bc5 ;
    mem[8'h40] <= 32'h9488f9e9 ;
    mem[8'h41] <= 32'hdbdf91f8 ;
    mem[8'h42] <= 32'ha2629cb ;
    mem[8'h43] <= 32'h457141da ;
    mem[8'h44] <= 32'had14441a ;
    mem[8'h45] <= 32'he2432c0b ;
    mem[8'h46] <= 32'h33ba9438 ;
    mem[8'h47] <= 32'h7cedfc29 ;
    mem[8'h48] <= 32'he7b1820f ;
    mem[8'h49] <= 32'ha8e6ea1e ;
    mem[8'h4a] <= 32'h791f522d ;
    mem[8'h4b] <= 32'h36483a3c ;
    mem[8'h4c] <= 32'hde2d3ffc ;
    mem[8'h4d] <= 32'h917a57ed ;
    mem[8'h4e] <= 32'h4083efde ;
    mem[8'h4f] <= 32'hfd487cf ;
    mem[8'h50] <= 32'h72fa0e25 ;
    mem[8'h51] <= 32'h3dad6634 ;
    mem[8'h52] <= 32'hec54de07 ;
    mem[8'h53] <= 32'ha303b616 ;
    mem[8'h54] <= 32'h4b66b3d6 ;
    mem[8'h55] <= 32'h431dbc7 ;
    mem[8'h56] <= 32'hd5c863f4 ;
    mem[8'h57] <= 32'h9a9f0be5 ;
    mem[8'h58] <= 32'h1c375c3 ;
    mem[8'h59] <= 32'h4e941dd2 ;
    mem[8'h5a] <= 32'h9f6da5e1 ;
    mem[8'h5b] <= 32'hd03acdf0 ;
    mem[8'h5c] <= 32'h385fc830 ;
    mem[8'h5d] <= 32'h7708a021 ;
    mem[8'h5e] <= 32'ha6f11812 ;
    mem[8'h5f] <= 32'he9a67003 ;
    mem[8'h60] <= 32'h5cac0bc6 ;
    mem[8'h61] <= 32'h13fb63d7 ;
    mem[8'h62] <= 32'hc202dbe4 ;
    mem[8'h63] <= 32'h8d55b3f5 ;
    mem[8'h64] <= 32'h6530b635 ;
    mem[8'h65] <= 32'h2a67de24 ;
    mem[8'h66] <= 32'hfb9e6617 ;
    mem[8'h67] <= 32'hb4c90e06 ;
    mem[8'h68] <= 32'h2f957020 ;
    mem[8'h69] <= 32'h60c21831 ;
    mem[8'h6a] <= 32'hb13ba002 ;
    mem[8'h6b] <= 32'hfe6cc813 ;
    mem[8'h6c] <= 32'h1609cdd3 ;
    mem[8'h6d] <= 32'h595ea5c2 ;
    mem[8'h6e] <= 32'h88a71df1 ;
    mem[8'h6f] <= 32'hc7f075e0 ;
    mem[8'h70] <= 32'hbadefc0a ;
    mem[8'h71] <= 32'hf589941b ;
    mem[8'h72] <= 32'h24702c28 ;
    mem[8'h73] <= 32'h6b274439 ;
    mem[8'h74] <= 32'h834241f9 ;
    mem[8'h75] <= 32'hcc1529e8 ;
    mem[8'h76] <= 32'h1dec91db ;
    mem[8'h77] <= 32'h52bbf9ca ;
    mem[8'h78] <= 32'hc9e787ec ;
    mem[8'h79] <= 32'h86b0effd ;
    mem[8'h7a] <= 32'h574957ce ;
    mem[8'h7b] <= 32'h181e3fdf ;
    mem[8'h7c] <= 32'hf07b3a1f ;
    mem[8'h7d] <= 32'hbf2c520e ;
    mem[8'h7e] <= 32'h6ed5ea3d ;
    mem[8'h7f] <= 32'h2182822c ;
    mem[8'h80] <= 32'h2dd0ee65 ;
    mem[8'h81] <= 32'h62878674 ;
    mem[8'h82] <= 32'hb37e3e47 ;
    mem[8'h83] <= 32'hfc295656 ;
    mem[8'h84] <= 32'h144c5396 ;
    mem[8'h85] <= 32'h5b1b3b87 ;
    mem[8'h86] <= 32'h8ae283b4 ;
    mem[8'h87] <= 32'hc5b5eba5 ;
    mem[8'h88] <= 32'h5ee99583 ;
    mem[8'h89] <= 32'h11befd92 ;
    mem[8'h8a] <= 32'hc04745a1 ;
    mem[8'h8b] <= 32'h8f102db0 ;
    mem[8'h8c] <= 32'h67752870 ;
    mem[8'h8d] <= 32'h28224061 ;
    mem[8'h8e] <= 32'hf9dbf852 ;
    mem[8'h8f] <= 32'hb68c9043 ;
    mem[8'h90] <= 32'hcba219a9 ;
    mem[8'h91] <= 32'h84f571b8 ;
    mem[8'h92] <= 32'h550cc98b ;
    mem[8'h93] <= 32'h1a5ba19a ;
    mem[8'h94] <= 32'hf23ea45a ;
    mem[8'h95] <= 32'hbd69cc4b ;
    mem[8'h96] <= 32'h6c907478 ;
    mem[8'h97] <= 32'h23c71c69 ;
    mem[8'h98] <= 32'hb89b624f ;
    mem[8'h99] <= 32'hf7cc0a5e ;
    mem[8'h9a] <= 32'h2635b26d ;
    mem[8'h9b] <= 32'h6962da7c ;
    mem[8'h9c] <= 32'h8107dfbc ;
    mem[8'h9d] <= 32'hce50b7ad ;
    mem[8'h9e] <= 32'h1fa90f9e ;
    mem[8'h9f] <= 32'h50fe678f ;
    mem[8'ha0] <= 32'he5f41c4a ;
    mem[8'ha1] <= 32'haaa3745b ;
    mem[8'ha2] <= 32'h7b5acc68 ;
    mem[8'ha3] <= 32'h340da479 ;
    mem[8'ha4] <= 32'hdc68a1b9 ;
    mem[8'ha5] <= 32'h933fc9a8 ;
    mem[8'ha6] <= 32'h42c6719b ;
    mem[8'ha7] <= 32'hd91198a ;
    mem[8'ha8] <= 32'h96cd67ac ;
    mem[8'ha9] <= 32'hd99a0fbd ;
    mem[8'haa] <= 32'h863b78e ;
    mem[8'hab] <= 32'h4734df9f ;
    mem[8'hac] <= 32'haf51da5f ;
    mem[8'had] <= 32'he006b24e ;
    mem[8'hae] <= 32'h31ff0a7d ;
    mem[8'haf] <= 32'h7ea8626c ;
    mem[8'hb0] <= 32'h386eb86 ;
    mem[8'hb1] <= 32'h4cd18397 ;
    mem[8'hb2] <= 32'h9d283ba4 ;
    mem[8'hb3] <= 32'hd27f53b5 ;
    mem[8'hb4] <= 32'h3a1a5675 ;
    mem[8'hb5] <= 32'h754d3e64 ;
    mem[8'hb6] <= 32'ha4b48657 ;
    mem[8'hb7] <= 32'hebe3ee46 ;
    mem[8'hb8] <= 32'h70bf9060 ;
    mem[8'hb9] <= 32'h3fe8f871 ;
    mem[8'hba] <= 32'hee114042 ;
    mem[8'hbb] <= 32'ha1462853 ;
    mem[8'hbc] <= 32'h49232d93 ;
    mem[8'hbd] <= 32'h6744582 ;
    mem[8'hbe] <= 32'hd78dfdb1 ;
    mem[8'hbf] <= 32'h98da95a0 ;
    mem[8'hc0] <= 32'hb958178c ;
    mem[8'hc1] <= 32'hf60f7f9d ;
    mem[8'hc2] <= 32'h27f6c7ae ;
    mem[8'hc3] <= 32'h68a1afbf ;
    mem[8'hc4] <= 32'h80c4aa7f ;
    mem[8'hc5] <= 32'hcf93c26e ;
    mem[8'hc6] <= 32'h1e6a7a5d ;
    mem[8'hc7] <= 32'h513d124c ;
    mem[8'hc8] <= 32'hca616c6a ;
    mem[8'hc9] <= 32'h8536047b ;
    mem[8'hca] <= 32'h54cfbc48 ;
    mem[8'hcb] <= 32'h1b98d459 ;
    mem[8'hcc] <= 32'hf3fdd199 ;
    mem[8'hcd] <= 32'hbcaab988 ;
    mem[8'hce] <= 32'h6d5301bb ;
    mem[8'hcf] <= 32'h220469aa ;
    mem[8'hd0] <= 32'h5f2ae040 ;
    mem[8'hd1] <= 32'h107d8851 ;
    mem[8'hd2] <= 32'hc1843062 ;
    mem[8'hd3] <= 32'h8ed35873 ;
    mem[8'hd4] <= 32'h66b65db3 ;
    mem[8'hd5] <= 32'h29e135a2 ;
    mem[8'hd6] <= 32'hf8188d91 ;
    mem[8'hd7] <= 32'hb74fe580 ;
    mem[8'hd8] <= 32'h2c139ba6 ;
    mem[8'hd9] <= 32'h6344f3b7 ;
    mem[8'hda] <= 32'hb2bd4b84 ;
    mem[8'hdb] <= 32'hfdea2395 ;
    mem[8'hdc] <= 32'h158f2655 ;
    mem[8'hdd] <= 32'h5ad84e44 ;
    mem[8'hde] <= 32'h8b21f677 ;
    mem[8'hdf] <= 32'hc4769e66 ;
    mem[8'he0] <= 32'h717ce5a3 ;
    mem[8'he1] <= 32'h3e2b8db2 ;
    mem[8'he2] <= 32'hefd23581 ;
    mem[8'he3] <= 32'ha0855d90 ;
    mem[8'he4] <= 32'h48e05850 ;
    mem[8'he5] <= 32'h7b73041 ;
    mem[8'he6] <= 32'hd64e8872 ;
    mem[8'he7] <= 32'h9919e063 ;
    mem[8'he8] <= 32'h2459e45 ;
    mem[8'he9] <= 32'h4d12f654 ;
    mem[8'hea] <= 32'h9ceb4e67 ;
    mem[8'heb] <= 32'hd3bc2676 ;
    mem[8'hec] <= 32'h3bd923b6 ;
    mem[8'hed] <= 32'h748e4ba7 ;
    mem[8'hee] <= 32'ha577f394 ;
    mem[8'hef] <= 32'hea209b85 ;
    mem[8'hf0] <= 32'h970e126f ;
    mem[8'hf1] <= 32'hd8597a7e ;
    mem[8'hf2] <= 32'h9a0c24d ;
    mem[8'hf3] <= 32'h46f7aa5c ;
    mem[8'hf4] <= 32'hae92af9c ;
    mem[8'hf5] <= 32'he1c5c78d ;
    mem[8'hf6] <= 32'h303c7fbe ;
    mem[8'hf7] <= 32'h7f6b17af ;
    mem[8'hf8] <= 32'he4376989 ;
    mem[8'hf9] <= 32'hab600198 ;
    mem[8'hfa] <= 32'h7a99b9ab ;
    mem[8'hfb] <= 32'h35ced1ba ;
    mem[8'hfc] <= 32'hddabd47a ;
    mem[8'hfd] <= 32'h92fcbc6b ;
    mem[8'hfe] <= 32'h43050458 ;
    mem[8'hff] <= 32'hc526c49 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
