module crctab_ev21
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'hf382b7f2 ;
    mem[8'h2] <= 32'he3c47253 ;
    mem[8'h3] <= 32'h1046c5a1 ;
    mem[8'h4] <= 32'hc349f911 ;
    mem[8'h5] <= 32'h30cb4ee3 ;
    mem[8'h6] <= 32'h208d8b42 ;
    mem[8'h7] <= 32'hd30f3cb0 ;
    mem[8'h8] <= 32'h8252ef95 ;
    mem[8'h9] <= 32'h71d05867 ;
    mem[8'ha] <= 32'h61969dc6 ;
    mem[8'hb] <= 32'h92142a34 ;
    mem[8'hc] <= 32'h411b1684 ;
    mem[8'hd] <= 32'hb299a176 ;
    mem[8'he] <= 32'ha2df64d7 ;
    mem[8'hf] <= 32'h515dd325 ;
    mem[8'h10] <= 32'h64c29d ;
    mem[8'h11] <= 32'hf3e6756f ;
    mem[8'h12] <= 32'he3a0b0ce ;
    mem[8'h13] <= 32'h1022073c ;
    mem[8'h14] <= 32'hc32d3b8c ;
    mem[8'h15] <= 32'h30af8c7e ;
    mem[8'h16] <= 32'h20e949df ;
    mem[8'h17] <= 32'hd36bfe2d ;
    mem[8'h18] <= 32'h82362d08 ;
    mem[8'h19] <= 32'h71b49afa ;
    mem[8'h1a] <= 32'h61f25f5b ;
    mem[8'h1b] <= 32'h9270e8a9 ;
    mem[8'h1c] <= 32'h417fd419 ;
    mem[8'h1d] <= 32'hb2fd63eb ;
    mem[8'h1e] <= 32'ha2bba64a ;
    mem[8'h1f] <= 32'h513911b8 ;
    mem[8'h20] <= 32'hc9853a ;
    mem[8'h21] <= 32'hf34b32c8 ;
    mem[8'h22] <= 32'he30df769 ;
    mem[8'h23] <= 32'h108f409b ;
    mem[8'h24] <= 32'hc3807c2b ;
    mem[8'h25] <= 32'h3002cbd9 ;
    mem[8'h26] <= 32'h20440e78 ;
    mem[8'h27] <= 32'hd3c6b98a ;
    mem[8'h28] <= 32'h829b6aaf ;
    mem[8'h29] <= 32'h7119dd5d ;
    mem[8'h2a] <= 32'h615f18fc ;
    mem[8'h2b] <= 32'h92ddaf0e ;
    mem[8'h2c] <= 32'h41d293be ;
    mem[8'h2d] <= 32'hb250244c ;
    mem[8'h2e] <= 32'ha216e1ed ;
    mem[8'h2f] <= 32'h5194561f ;
    mem[8'h30] <= 32'had47a7 ;
    mem[8'h31] <= 32'hf32ff055 ;
    mem[8'h32] <= 32'he36935f4 ;
    mem[8'h33] <= 32'h10eb8206 ;
    mem[8'h34] <= 32'hc3e4beb6 ;
    mem[8'h35] <= 32'h30660944 ;
    mem[8'h36] <= 32'h2020cce5 ;
    mem[8'h37] <= 32'hd3a27b17 ;
    mem[8'h38] <= 32'h82ffa832 ;
    mem[8'h39] <= 32'h717d1fc0 ;
    mem[8'h3a] <= 32'h613bda61 ;
    mem[8'h3b] <= 32'h92b96d93 ;
    mem[8'h3c] <= 32'h41b65123 ;
    mem[8'h3d] <= 32'hb234e6d1 ;
    mem[8'h3e] <= 32'ha2722370 ;
    mem[8'h3f] <= 32'h51f09482 ;
    mem[8'h40] <= 32'h1930a74 ;
    mem[8'h41] <= 32'hf211bd86 ;
    mem[8'h42] <= 32'he2577827 ;
    mem[8'h43] <= 32'h11d5cfd5 ;
    mem[8'h44] <= 32'hc2daf365 ;
    mem[8'h45] <= 32'h31584497 ;
    mem[8'h46] <= 32'h211e8136 ;
    mem[8'h47] <= 32'hd29c36c4 ;
    mem[8'h48] <= 32'h83c1e5e1 ;
    mem[8'h49] <= 32'h70435213 ;
    mem[8'h4a] <= 32'h600597b2 ;
    mem[8'h4b] <= 32'h93872040 ;
    mem[8'h4c] <= 32'h40881cf0 ;
    mem[8'h4d] <= 32'hb30aab02 ;
    mem[8'h4e] <= 32'ha34c6ea3 ;
    mem[8'h4f] <= 32'h50ced951 ;
    mem[8'h50] <= 32'h1f7c8e9 ;
    mem[8'h51] <= 32'hf2757f1b ;
    mem[8'h52] <= 32'he233baba ;
    mem[8'h53] <= 32'h11b10d48 ;
    mem[8'h54] <= 32'hc2be31f8 ;
    mem[8'h55] <= 32'h313c860a ;
    mem[8'h56] <= 32'h217a43ab ;
    mem[8'h57] <= 32'hd2f8f459 ;
    mem[8'h58] <= 32'h83a5277c ;
    mem[8'h59] <= 32'h7027908e ;
    mem[8'h5a] <= 32'h6061552f ;
    mem[8'h5b] <= 32'h93e3e2dd ;
    mem[8'h5c] <= 32'h40ecde6d ;
    mem[8'h5d] <= 32'hb36e699f ;
    mem[8'h5e] <= 32'ha328ac3e ;
    mem[8'h5f] <= 32'h50aa1bcc ;
    mem[8'h60] <= 32'h15a8f4e ;
    mem[8'h61] <= 32'hf2d838bc ;
    mem[8'h62] <= 32'he29efd1d ;
    mem[8'h63] <= 32'h111c4aef ;
    mem[8'h64] <= 32'hc213765f ;
    mem[8'h65] <= 32'h3191c1ad ;
    mem[8'h66] <= 32'h21d7040c ;
    mem[8'h67] <= 32'hd255b3fe ;
    mem[8'h68] <= 32'h830860db ;
    mem[8'h69] <= 32'h708ad729 ;
    mem[8'h6a] <= 32'h60cc1288 ;
    mem[8'h6b] <= 32'h934ea57a ;
    mem[8'h6c] <= 32'h404199ca ;
    mem[8'h6d] <= 32'hb3c32e38 ;
    mem[8'h6e] <= 32'ha385eb99 ;
    mem[8'h6f] <= 32'h50075c6b ;
    mem[8'h70] <= 32'h13e4dd3 ;
    mem[8'h71] <= 32'hf2bcfa21 ;
    mem[8'h72] <= 32'he2fa3f80 ;
    mem[8'h73] <= 32'h11788872 ;
    mem[8'h74] <= 32'hc277b4c2 ;
    mem[8'h75] <= 32'h31f50330 ;
    mem[8'h76] <= 32'h21b3c691 ;
    mem[8'h77] <= 32'hd2317163 ;
    mem[8'h78] <= 32'h836ca246 ;
    mem[8'h79] <= 32'h70ee15b4 ;
    mem[8'h7a] <= 32'h60a8d015 ;
    mem[8'h7b] <= 32'h932a67e7 ;
    mem[8'h7c] <= 32'h40255b57 ;
    mem[8'h7d] <= 32'hb3a7eca5 ;
    mem[8'h7e] <= 32'ha3e12904 ;
    mem[8'h7f] <= 32'h50639ef6 ;
    mem[8'h80] <= 32'h32614e8 ;
    mem[8'h81] <= 32'hf0a4a31a ;
    mem[8'h82] <= 32'he0e266bb ;
    mem[8'h83] <= 32'h1360d149 ;
    mem[8'h84] <= 32'hc06fedf9 ;
    mem[8'h85] <= 32'h33ed5a0b ;
    mem[8'h86] <= 32'h23ab9faa ;
    mem[8'h87] <= 32'hd0292858 ;
    mem[8'h88] <= 32'h8174fb7d ;
    mem[8'h89] <= 32'h72f64c8f ;
    mem[8'h8a] <= 32'h62b0892e ;
    mem[8'h8b] <= 32'h91323edc ;
    mem[8'h8c] <= 32'h423d026c ;
    mem[8'h8d] <= 32'hb1bfb59e ;
    mem[8'h8e] <= 32'ha1f9703f ;
    mem[8'h8f] <= 32'h527bc7cd ;
    mem[8'h90] <= 32'h342d675 ;
    mem[8'h91] <= 32'hf0c06187 ;
    mem[8'h92] <= 32'he086a426 ;
    mem[8'h93] <= 32'h130413d4 ;
    mem[8'h94] <= 32'hc00b2f64 ;
    mem[8'h95] <= 32'h33899896 ;
    mem[8'h96] <= 32'h23cf5d37 ;
    mem[8'h97] <= 32'hd04deac5 ;
    mem[8'h98] <= 32'h811039e0 ;
    mem[8'h99] <= 32'h72928e12 ;
    mem[8'h9a] <= 32'h62d44bb3 ;
    mem[8'h9b] <= 32'h9156fc41 ;
    mem[8'h9c] <= 32'h4259c0f1 ;
    mem[8'h9d] <= 32'hb1db7703 ;
    mem[8'h9e] <= 32'ha19db2a2 ;
    mem[8'h9f] <= 32'h521f0550 ;
    mem[8'ha0] <= 32'h3ef91d2 ;
    mem[8'ha1] <= 32'hf06d2620 ;
    mem[8'ha2] <= 32'he02be381 ;
    mem[8'ha3] <= 32'h13a95473 ;
    mem[8'ha4] <= 32'hc0a668c3 ;
    mem[8'ha5] <= 32'h3324df31 ;
    mem[8'ha6] <= 32'h23621a90 ;
    mem[8'ha7] <= 32'hd0e0ad62 ;
    mem[8'ha8] <= 32'h81bd7e47 ;
    mem[8'ha9] <= 32'h723fc9b5 ;
    mem[8'haa] <= 32'h62790c14 ;
    mem[8'hab] <= 32'h91fbbbe6 ;
    mem[8'hac] <= 32'h42f48756 ;
    mem[8'had] <= 32'hb17630a4 ;
    mem[8'hae] <= 32'ha130f505 ;
    mem[8'haf] <= 32'h52b242f7 ;
    mem[8'hb0] <= 32'h38b534f ;
    mem[8'hb1] <= 32'hf009e4bd ;
    mem[8'hb2] <= 32'he04f211c ;
    mem[8'hb3] <= 32'h13cd96ee ;
    mem[8'hb4] <= 32'hc0c2aa5e ;
    mem[8'hb5] <= 32'h33401dac ;
    mem[8'hb6] <= 32'h2306d80d ;
    mem[8'hb7] <= 32'hd0846fff ;
    mem[8'hb8] <= 32'h81d9bcda ;
    mem[8'hb9] <= 32'h725b0b28 ;
    mem[8'hba] <= 32'h621dce89 ;
    mem[8'hbb] <= 32'h919f797b ;
    mem[8'hbc] <= 32'h429045cb ;
    mem[8'hbd] <= 32'hb112f239 ;
    mem[8'hbe] <= 32'ha1543798 ;
    mem[8'hbf] <= 32'h52d6806a ;
    mem[8'hc0] <= 32'h2b51e9c ;
    mem[8'hc1] <= 32'hf137a96e ;
    mem[8'hc2] <= 32'he1716ccf ;
    mem[8'hc3] <= 32'h12f3db3d ;
    mem[8'hc4] <= 32'hc1fce78d ;
    mem[8'hc5] <= 32'h327e507f ;
    mem[8'hc6] <= 32'h223895de ;
    mem[8'hc7] <= 32'hd1ba222c ;
    mem[8'hc8] <= 32'h80e7f109 ;
    mem[8'hc9] <= 32'h736546fb ;
    mem[8'hca] <= 32'h6323835a ;
    mem[8'hcb] <= 32'h90a134a8 ;
    mem[8'hcc] <= 32'h43ae0818 ;
    mem[8'hcd] <= 32'hb02cbfea ;
    mem[8'hce] <= 32'ha06a7a4b ;
    mem[8'hcf] <= 32'h53e8cdb9 ;
    mem[8'hd0] <= 32'h2d1dc01 ;
    mem[8'hd1] <= 32'hf1536bf3 ;
    mem[8'hd2] <= 32'he115ae52 ;
    mem[8'hd3] <= 32'h129719a0 ;
    mem[8'hd4] <= 32'hc1982510 ;
    mem[8'hd5] <= 32'h321a92e2 ;
    mem[8'hd6] <= 32'h225c5743 ;
    mem[8'hd7] <= 32'hd1dee0b1 ;
    mem[8'hd8] <= 32'h80833394 ;
    mem[8'hd9] <= 32'h73018466 ;
    mem[8'hda] <= 32'h634741c7 ;
    mem[8'hdb] <= 32'h90c5f635 ;
    mem[8'hdc] <= 32'h43caca85 ;
    mem[8'hdd] <= 32'hb0487d77 ;
    mem[8'hde] <= 32'ha00eb8d6 ;
    mem[8'hdf] <= 32'h538c0f24 ;
    mem[8'he0] <= 32'h27c9ba6 ;
    mem[8'he1] <= 32'hf1fe2c54 ;
    mem[8'he2] <= 32'he1b8e9f5 ;
    mem[8'he3] <= 32'h123a5e07 ;
    mem[8'he4] <= 32'hc13562b7 ;
    mem[8'he5] <= 32'h32b7d545 ;
    mem[8'he6] <= 32'h22f110e4 ;
    mem[8'he7] <= 32'hd173a716 ;
    mem[8'he8] <= 32'h802e7433 ;
    mem[8'he9] <= 32'h73acc3c1 ;
    mem[8'hea] <= 32'h63ea0660 ;
    mem[8'heb] <= 32'h9068b192 ;
    mem[8'hec] <= 32'h43678d22 ;
    mem[8'hed] <= 32'hb0e53ad0 ;
    mem[8'hee] <= 32'ha0a3ff71 ;
    mem[8'hef] <= 32'h53214883 ;
    mem[8'hf0] <= 32'h218593b ;
    mem[8'hf1] <= 32'hf19aeec9 ;
    mem[8'hf2] <= 32'he1dc2b68 ;
    mem[8'hf3] <= 32'h125e9c9a ;
    mem[8'hf4] <= 32'hc151a02a ;
    mem[8'hf5] <= 32'h32d317d8 ;
    mem[8'hf6] <= 32'h2295d279 ;
    mem[8'hf7] <= 32'hd117658b ;
    mem[8'hf8] <= 32'h804ab6ae ;
    mem[8'hf9] <= 32'h73c8015c ;
    mem[8'hfa] <= 32'h638ec4fd ;
    mem[8'hfb] <= 32'h900c730f ;
    mem[8'hfc] <= 32'h43034fbf ;
    mem[8'hfd] <= 32'hb081f84d ;
    mem[8'hfe] <= 32'ha0c73dec ;
    mem[8'hff] <= 32'h53458a1e ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
