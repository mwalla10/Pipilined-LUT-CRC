module crctab_ev8
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'hf200aa66 ;
    mem[8'h2] <= 32'he0c0497b ;
    mem[8'h3] <= 32'h12c0e31d ;
    mem[8'h4] <= 32'hc5418f41 ;
    mem[8'h5] <= 32'h37412527 ;
    mem[8'h6] <= 32'h2581c63a ;
    mem[8'h7] <= 32'hd7816c5c ;
    mem[8'h8] <= 32'h8e420335 ;
    mem[8'h9] <= 32'h7c42a953 ;
    mem[8'ha] <= 32'h6e824a4e ;
    mem[8'hb] <= 32'h9c82e028 ;
    mem[8'hc] <= 32'h4b038c74 ;
    mem[8'hd] <= 32'hb9032612 ;
    mem[8'he] <= 32'habc3c50f ;
    mem[8'hf] <= 32'h59c36f69 ;
    mem[8'h10] <= 32'h18451bdd ;
    mem[8'h11] <= 32'hea45b1bb ;
    mem[8'h12] <= 32'hf88552a6 ;
    mem[8'h13] <= 32'ha85f8c0 ;
    mem[8'h14] <= 32'hdd04949c ;
    mem[8'h15] <= 32'h2f043efa ;
    mem[8'h16] <= 32'h3dc4dde7 ;
    mem[8'h17] <= 32'hcfc47781 ;
    mem[8'h18] <= 32'h960718e8 ;
    mem[8'h19] <= 32'h6407b28e ;
    mem[8'h1a] <= 32'h76c75193 ;
    mem[8'h1b] <= 32'h84c7fbf5 ;
    mem[8'h1c] <= 32'h534697a9 ;
    mem[8'h1d] <= 32'ha1463dcf ;
    mem[8'h1e] <= 32'hb386ded2 ;
    mem[8'h1f] <= 32'h418674b4 ;
    mem[8'h20] <= 32'h308a37ba ;
    mem[8'h21] <= 32'hc28a9ddc ;
    mem[8'h22] <= 32'hd04a7ec1 ;
    mem[8'h23] <= 32'h224ad4a7 ;
    mem[8'h24] <= 32'hf5cbb8fb ;
    mem[8'h25] <= 32'h7cb129d ;
    mem[8'h26] <= 32'h150bf180 ;
    mem[8'h27] <= 32'he70b5be6 ;
    mem[8'h28] <= 32'hbec8348f ;
    mem[8'h29] <= 32'h4cc89ee9 ;
    mem[8'h2a] <= 32'h5e087df4 ;
    mem[8'h2b] <= 32'hac08d792 ;
    mem[8'h2c] <= 32'h7b89bbce ;
    mem[8'h2d] <= 32'h898911a8 ;
    mem[8'h2e] <= 32'h9b49f2b5 ;
    mem[8'h2f] <= 32'h694958d3 ;
    mem[8'h30] <= 32'h28cf2c67 ;
    mem[8'h31] <= 32'hdacf8601 ;
    mem[8'h32] <= 32'hc80f651c ;
    mem[8'h33] <= 32'h3a0fcf7a ;
    mem[8'h34] <= 32'hed8ea326 ;
    mem[8'h35] <= 32'h1f8e0940 ;
    mem[8'h36] <= 32'hd4eea5d ;
    mem[8'h37] <= 32'hff4e403b ;
    mem[8'h38] <= 32'ha68d2f52 ;
    mem[8'h39] <= 32'h548d8534 ;
    mem[8'h3a] <= 32'h464d6629 ;
    mem[8'h3b] <= 32'hb44dcc4f ;
    mem[8'h3c] <= 32'h63cca013 ;
    mem[8'h3d] <= 32'h91cc0a75 ;
    mem[8'h3e] <= 32'h830ce968 ;
    mem[8'h3f] <= 32'h710c430e ;
    mem[8'h40] <= 32'h61146f74 ;
    mem[8'h41] <= 32'h9314c512 ;
    mem[8'h42] <= 32'h81d4260f ;
    mem[8'h43] <= 32'h73d48c69 ;
    mem[8'h44] <= 32'ha455e035 ;
    mem[8'h45] <= 32'h56554a53 ;
    mem[8'h46] <= 32'h4495a94e ;
    mem[8'h47] <= 32'hb6950328 ;
    mem[8'h48] <= 32'hef566c41 ;
    mem[8'h49] <= 32'h1d56c627 ;
    mem[8'h4a] <= 32'hf96253a ;
    mem[8'h4b] <= 32'hfd968f5c ;
    mem[8'h4c] <= 32'h2a17e300 ;
    mem[8'h4d] <= 32'hd8174966 ;
    mem[8'h4e] <= 32'hcad7aa7b ;
    mem[8'h4f] <= 32'h38d7001d ;
    mem[8'h50] <= 32'h795174a9 ;
    mem[8'h51] <= 32'h8b51decf ;
    mem[8'h52] <= 32'h99913dd2 ;
    mem[8'h53] <= 32'h6b9197b4 ;
    mem[8'h54] <= 32'hbc10fbe8 ;
    mem[8'h55] <= 32'h4e10518e ;
    mem[8'h56] <= 32'h5cd0b293 ;
    mem[8'h57] <= 32'haed018f5 ;
    mem[8'h58] <= 32'hf713779c ;
    mem[8'h59] <= 32'h513ddfa ;
    mem[8'h5a] <= 32'h17d33ee7 ;
    mem[8'h5b] <= 32'he5d39481 ;
    mem[8'h5c] <= 32'h3252f8dd ;
    mem[8'h5d] <= 32'hc05252bb ;
    mem[8'h5e] <= 32'hd292b1a6 ;
    mem[8'h5f] <= 32'h20921bc0 ;
    mem[8'h60] <= 32'h519e58ce ;
    mem[8'h61] <= 32'ha39ef2a8 ;
    mem[8'h62] <= 32'hb15e11b5 ;
    mem[8'h63] <= 32'h435ebbd3 ;
    mem[8'h64] <= 32'h94dfd78f ;
    mem[8'h65] <= 32'h66df7de9 ;
    mem[8'h66] <= 32'h741f9ef4 ;
    mem[8'h67] <= 32'h861f3492 ;
    mem[8'h68] <= 32'hdfdc5bfb ;
    mem[8'h69] <= 32'h2ddcf19d ;
    mem[8'h6a] <= 32'h3f1c1280 ;
    mem[8'h6b] <= 32'hcd1cb8e6 ;
    mem[8'h6c] <= 32'h1a9dd4ba ;
    mem[8'h6d] <= 32'he89d7edc ;
    mem[8'h6e] <= 32'hfa5d9dc1 ;
    mem[8'h6f] <= 32'h85d37a7 ;
    mem[8'h70] <= 32'h49db4313 ;
    mem[8'h71] <= 32'hbbdbe975 ;
    mem[8'h72] <= 32'ha91b0a68 ;
    mem[8'h73] <= 32'h5b1ba00e ;
    mem[8'h74] <= 32'h8c9acc52 ;
    mem[8'h75] <= 32'h7e9a6634 ;
    mem[8'h76] <= 32'h6c5a8529 ;
    mem[8'h77] <= 32'h9e5a2f4f ;
    mem[8'h78] <= 32'hc7994026 ;
    mem[8'h79] <= 32'h3599ea40 ;
    mem[8'h7a] <= 32'h2759095d ;
    mem[8'h7b] <= 32'hd559a33b ;
    mem[8'h7c] <= 32'h2d8cf67 ;
    mem[8'h7d] <= 32'hf0d86501 ;
    mem[8'h7e] <= 32'he218861c ;
    mem[8'h7f] <= 32'h10182c7a ;
    mem[8'h80] <= 32'hc228dee8 ;
    mem[8'h81] <= 32'h3028748e ;
    mem[8'h82] <= 32'h22e89793 ;
    mem[8'h83] <= 32'hd0e83df5 ;
    mem[8'h84] <= 32'h76951a9 ;
    mem[8'h85] <= 32'hf569fbcf ;
    mem[8'h86] <= 32'he7a918d2 ;
    mem[8'h87] <= 32'h15a9b2b4 ;
    mem[8'h88] <= 32'h4c6adddd ;
    mem[8'h89] <= 32'hbe6a77bb ;
    mem[8'h8a] <= 32'hacaa94a6 ;
    mem[8'h8b] <= 32'h5eaa3ec0 ;
    mem[8'h8c] <= 32'h892b529c ;
    mem[8'h8d] <= 32'h7b2bf8fa ;
    mem[8'h8e] <= 32'h69eb1be7 ;
    mem[8'h8f] <= 32'h9bebb181 ;
    mem[8'h90] <= 32'hda6dc535 ;
    mem[8'h91] <= 32'h286d6f53 ;
    mem[8'h92] <= 32'h3aad8c4e ;
    mem[8'h93] <= 32'hc8ad2628 ;
    mem[8'h94] <= 32'h1f2c4a74 ;
    mem[8'h95] <= 32'hed2ce012 ;
    mem[8'h96] <= 32'hffec030f ;
    mem[8'h97] <= 32'hdeca969 ;
    mem[8'h98] <= 32'h542fc600 ;
    mem[8'h99] <= 32'ha62f6c66 ;
    mem[8'h9a] <= 32'hb4ef8f7b ;
    mem[8'h9b] <= 32'h46ef251d ;
    mem[8'h9c] <= 32'h916e4941 ;
    mem[8'h9d] <= 32'h636ee327 ;
    mem[8'h9e] <= 32'h71ae003a ;
    mem[8'h9f] <= 32'h83aeaa5c ;
    mem[8'ha0] <= 32'hf2a2e952 ;
    mem[8'ha1] <= 32'ha24334 ;
    mem[8'ha2] <= 32'h1262a029 ;
    mem[8'ha3] <= 32'he0620a4f ;
    mem[8'ha4] <= 32'h37e36613 ;
    mem[8'ha5] <= 32'hc5e3cc75 ;
    mem[8'ha6] <= 32'hd7232f68 ;
    mem[8'ha7] <= 32'h2523850e ;
    mem[8'ha8] <= 32'h7ce0ea67 ;
    mem[8'ha9] <= 32'h8ee04001 ;
    mem[8'haa] <= 32'h9c20a31c ;
    mem[8'hab] <= 32'h6e20097a ;
    mem[8'hac] <= 32'hb9a16526 ;
    mem[8'had] <= 32'h4ba1cf40 ;
    mem[8'hae] <= 32'h59612c5d ;
    mem[8'haf] <= 32'hab61863b ;
    mem[8'hb0] <= 32'heae7f28f ;
    mem[8'hb1] <= 32'h18e758e9 ;
    mem[8'hb2] <= 32'ha27bbf4 ;
    mem[8'hb3] <= 32'hf8271192 ;
    mem[8'hb4] <= 32'h2fa67dce ;
    mem[8'hb5] <= 32'hdda6d7a8 ;
    mem[8'hb6] <= 32'hcf6634b5 ;
    mem[8'hb7] <= 32'h3d669ed3 ;
    mem[8'hb8] <= 32'h64a5f1ba ;
    mem[8'hb9] <= 32'h96a55bdc ;
    mem[8'hba] <= 32'h8465b8c1 ;
    mem[8'hbb] <= 32'h766512a7 ;
    mem[8'hbc] <= 32'ha1e47efb ;
    mem[8'hbd] <= 32'h53e4d49d ;
    mem[8'hbe] <= 32'h41243780 ;
    mem[8'hbf] <= 32'hb3249de6 ;
    mem[8'hc0] <= 32'ha33cb19c ;
    mem[8'hc1] <= 32'h513c1bfa ;
    mem[8'hc2] <= 32'h43fcf8e7 ;
    mem[8'hc3] <= 32'hb1fc5281 ;
    mem[8'hc4] <= 32'h667d3edd ;
    mem[8'hc5] <= 32'h947d94bb ;
    mem[8'hc6] <= 32'h86bd77a6 ;
    mem[8'hc7] <= 32'h74bdddc0 ;
    mem[8'hc8] <= 32'h2d7eb2a9 ;
    mem[8'hc9] <= 32'hdf7e18cf ;
    mem[8'hca] <= 32'hcdbefbd2 ;
    mem[8'hcb] <= 32'h3fbe51b4 ;
    mem[8'hcc] <= 32'he83f3de8 ;
    mem[8'hcd] <= 32'h1a3f978e ;
    mem[8'hce] <= 32'h8ff7493 ;
    mem[8'hcf] <= 32'hfaffdef5 ;
    mem[8'hd0] <= 32'hbb79aa41 ;
    mem[8'hd1] <= 32'h49790027 ;
    mem[8'hd2] <= 32'h5bb9e33a ;
    mem[8'hd3] <= 32'ha9b9495c ;
    mem[8'hd4] <= 32'h7e382500 ;
    mem[8'hd5] <= 32'h8c388f66 ;
    mem[8'hd6] <= 32'h9ef86c7b ;
    mem[8'hd7] <= 32'h6cf8c61d ;
    mem[8'hd8] <= 32'h353ba974 ;
    mem[8'hd9] <= 32'hc73b0312 ;
    mem[8'hda] <= 32'hd5fbe00f ;
    mem[8'hdb] <= 32'h27fb4a69 ;
    mem[8'hdc] <= 32'hf07a2635 ;
    mem[8'hdd] <= 32'h27a8c53 ;
    mem[8'hde] <= 32'h10ba6f4e ;
    mem[8'hdf] <= 32'he2bac528 ;
    mem[8'he0] <= 32'h93b68626 ;
    mem[8'he1] <= 32'h61b62c40 ;
    mem[8'he2] <= 32'h7376cf5d ;
    mem[8'he3] <= 32'h8176653b ;
    mem[8'he4] <= 32'h56f70967 ;
    mem[8'he5] <= 32'ha4f7a301 ;
    mem[8'he6] <= 32'hb637401c ;
    mem[8'he7] <= 32'h4437ea7a ;
    mem[8'he8] <= 32'h1df48513 ;
    mem[8'he9] <= 32'heff42f75 ;
    mem[8'hea] <= 32'hfd34cc68 ;
    mem[8'heb] <= 32'hf34660e ;
    mem[8'hec] <= 32'hd8b50a52 ;
    mem[8'hed] <= 32'h2ab5a034 ;
    mem[8'hee] <= 32'h38754329 ;
    mem[8'hef] <= 32'hca75e94f ;
    mem[8'hf0] <= 32'h8bf39dfb ;
    mem[8'hf1] <= 32'h79f3379d ;
    mem[8'hf2] <= 32'h6b33d480 ;
    mem[8'hf3] <= 32'h99337ee6 ;
    mem[8'hf4] <= 32'h4eb212ba ;
    mem[8'hf5] <= 32'hbcb2b8dc ;
    mem[8'hf6] <= 32'hae725bc1 ;
    mem[8'hf7] <= 32'h5c72f1a7 ;
    mem[8'hf8] <= 32'h5b19ece ;
    mem[8'hf9] <= 32'hf7b134a8 ;
    mem[8'hfa] <= 32'he571d7b5 ;
    mem[8'hfb] <= 32'h17717dd3 ;
    mem[8'hfc] <= 32'hc0f0118f ;
    mem[8'hfd] <= 32'h32f0bbe9 ;
    mem[8'hfe] <= 32'h203058f4 ;
    mem[8'hff] <= 32'hd230f292 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
