module crctab_ev28
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h75be46b7 ;
    mem[8'h2] <= 32'heb7c8d6e ;
    mem[8'h3] <= 32'h9ec2cbd9 ;
    mem[8'h4] <= 32'hd238076b ;
    mem[8'h5] <= 32'ha78641dc ;
    mem[8'h6] <= 32'h39448a05 ;
    mem[8'h7] <= 32'h4cfaccb2 ;
    mem[8'h8] <= 32'ha0b11361 ;
    mem[8'h9] <= 32'hd50f55d6 ;
    mem[8'ha] <= 32'h4bcd9e0f ;
    mem[8'hb] <= 32'h3e73d8b8 ;
    mem[8'hc] <= 32'h7289140a ;
    mem[8'hd] <= 32'h73752bd ;
    mem[8'he] <= 32'h99f59964 ;
    mem[8'hf] <= 32'hec4bdfd3 ;
    mem[8'h10] <= 32'h45a33b75 ;
    mem[8'h11] <= 32'h301d7dc2 ;
    mem[8'h12] <= 32'haedfb61b ;
    mem[8'h13] <= 32'hdb61f0ac ;
    mem[8'h14] <= 32'h979b3c1e ;
    mem[8'h15] <= 32'he2257aa9 ;
    mem[8'h16] <= 32'h7ce7b170 ;
    mem[8'h17] <= 32'h959f7c7 ;
    mem[8'h18] <= 32'he5122814 ;
    mem[8'h19] <= 32'h90ac6ea3 ;
    mem[8'h1a] <= 32'he6ea57a ;
    mem[8'h1b] <= 32'h7bd0e3cd ;
    mem[8'h1c] <= 32'h372a2f7f ;
    mem[8'h1d] <= 32'h429469c8 ;
    mem[8'h1e] <= 32'hdc56a211 ;
    mem[8'h1f] <= 32'ha9e8e4a6 ;
    mem[8'h20] <= 32'h8b4676ea ;
    mem[8'h21] <= 32'hfef8305d ;
    mem[8'h22] <= 32'h603afb84 ;
    mem[8'h23] <= 32'h1584bd33 ;
    mem[8'h24] <= 32'h597e7181 ;
    mem[8'h25] <= 32'h2cc03736 ;
    mem[8'h26] <= 32'hb202fcef ;
    mem[8'h27] <= 32'hc7bcba58 ;
    mem[8'h28] <= 32'h2bf7658b ;
    mem[8'h29] <= 32'h5e49233c ;
    mem[8'h2a] <= 32'hc08be8e5 ;
    mem[8'h2b] <= 32'hb535ae52 ;
    mem[8'h2c] <= 32'hf9cf62e0 ;
    mem[8'h2d] <= 32'h8c712457 ;
    mem[8'h2e] <= 32'h12b3ef8e ;
    mem[8'h2f] <= 32'h670da939 ;
    mem[8'h30] <= 32'hcee54d9f ;
    mem[8'h31] <= 32'hbb5b0b28 ;
    mem[8'h32] <= 32'h2599c0f1 ;
    mem[8'h33] <= 32'h50278646 ;
    mem[8'h34] <= 32'h1cdd4af4 ;
    mem[8'h35] <= 32'h69630c43 ;
    mem[8'h36] <= 32'hf7a1c79a ;
    mem[8'h37] <= 32'h821f812d ;
    mem[8'h38] <= 32'h6e545efe ;
    mem[8'h39] <= 32'h1bea1849 ;
    mem[8'h3a] <= 32'h8528d390 ;
    mem[8'h3b] <= 32'hf0969527 ;
    mem[8'h3c] <= 32'hbc6c5995 ;
    mem[8'h3d] <= 32'hc9d21f22 ;
    mem[8'h3e] <= 32'h5710d4fb ;
    mem[8'h3f] <= 32'h22ae924c ;
    mem[8'h40] <= 32'h124df063 ;
    mem[8'h41] <= 32'h67f3b6d4 ;
    mem[8'h42] <= 32'hf9317d0d ;
    mem[8'h43] <= 32'h8c8f3bba ;
    mem[8'h44] <= 32'hc075f708 ;
    mem[8'h45] <= 32'hb5cbb1bf ;
    mem[8'h46] <= 32'h2b097a66 ;
    mem[8'h47] <= 32'h5eb73cd1 ;
    mem[8'h48] <= 32'hb2fce302 ;
    mem[8'h49] <= 32'hc742a5b5 ;
    mem[8'h4a] <= 32'h59806e6c ;
    mem[8'h4b] <= 32'h2c3e28db ;
    mem[8'h4c] <= 32'h60c4e469 ;
    mem[8'h4d] <= 32'h157aa2de ;
    mem[8'h4e] <= 32'h8bb86907 ;
    mem[8'h4f] <= 32'hfe062fb0 ;
    mem[8'h50] <= 32'h57eecb16 ;
    mem[8'h51] <= 32'h22508da1 ;
    mem[8'h52] <= 32'hbc924678 ;
    mem[8'h53] <= 32'hc92c00cf ;
    mem[8'h54] <= 32'h85d6cc7d ;
    mem[8'h55] <= 32'hf0688aca ;
    mem[8'h56] <= 32'h6eaa4113 ;
    mem[8'h57] <= 32'h1b1407a4 ;
    mem[8'h58] <= 32'hf75fd877 ;
    mem[8'h59] <= 32'h82e19ec0 ;
    mem[8'h5a] <= 32'h1c235519 ;
    mem[8'h5b] <= 32'h699d13ae ;
    mem[8'h5c] <= 32'h2567df1c ;
    mem[8'h5d] <= 32'h50d999ab ;
    mem[8'h5e] <= 32'hce1b5272 ;
    mem[8'h5f] <= 32'hbba514c5 ;
    mem[8'h60] <= 32'h990b8689 ;
    mem[8'h61] <= 32'hecb5c03e ;
    mem[8'h62] <= 32'h72770be7 ;
    mem[8'h63] <= 32'h7c94d50 ;
    mem[8'h64] <= 32'h4b3381e2 ;
    mem[8'h65] <= 32'h3e8dc755 ;
    mem[8'h66] <= 32'ha04f0c8c ;
    mem[8'h67] <= 32'hd5f14a3b ;
    mem[8'h68] <= 32'h39ba95e8 ;
    mem[8'h69] <= 32'h4c04d35f ;
    mem[8'h6a] <= 32'hd2c61886 ;
    mem[8'h6b] <= 32'ha7785e31 ;
    mem[8'h6c] <= 32'heb829283 ;
    mem[8'h6d] <= 32'h9e3cd434 ;
    mem[8'h6e] <= 32'hfe1fed ;
    mem[8'h6f] <= 32'h7540595a ;
    mem[8'h70] <= 32'hdca8bdfc ;
    mem[8'h71] <= 32'ha916fb4b ;
    mem[8'h72] <= 32'h37d43092 ;
    mem[8'h73] <= 32'h426a7625 ;
    mem[8'h74] <= 32'he90ba97 ;
    mem[8'h75] <= 32'h7b2efc20 ;
    mem[8'h76] <= 32'he5ec37f9 ;
    mem[8'h77] <= 32'h9052714e ;
    mem[8'h78] <= 32'h7c19ae9d ;
    mem[8'h79] <= 32'h9a7e82a ;
    mem[8'h7a] <= 32'h976523f3 ;
    mem[8'h7b] <= 32'he2db6544 ;
    mem[8'h7c] <= 32'hae21a9f6 ;
    mem[8'h7d] <= 32'hdb9fef41 ;
    mem[8'h7e] <= 32'h455d2498 ;
    mem[8'h7f] <= 32'h30e3622f ;
    mem[8'h80] <= 32'h249be0c6 ;
    mem[8'h81] <= 32'h5125a671 ;
    mem[8'h82] <= 32'hcfe76da8 ;
    mem[8'h83] <= 32'hba592b1f ;
    mem[8'h84] <= 32'hf6a3e7ad ;
    mem[8'h85] <= 32'h831da11a ;
    mem[8'h86] <= 32'h1ddf6ac3 ;
    mem[8'h87] <= 32'h68612c74 ;
    mem[8'h88] <= 32'h842af3a7 ;
    mem[8'h89] <= 32'hf194b510 ;
    mem[8'h8a] <= 32'h6f567ec9 ;
    mem[8'h8b] <= 32'h1ae8387e ;
    mem[8'h8c] <= 32'h5612f4cc ;
    mem[8'h8d] <= 32'h23acb27b ;
    mem[8'h8e] <= 32'hbd6e79a2 ;
    mem[8'h8f] <= 32'hc8d03f15 ;
    mem[8'h90] <= 32'h6138dbb3 ;
    mem[8'h91] <= 32'h14869d04 ;
    mem[8'h92] <= 32'h8a4456dd ;
    mem[8'h93] <= 32'hfffa106a ;
    mem[8'h94] <= 32'hb300dcd8 ;
    mem[8'h95] <= 32'hc6be9a6f ;
    mem[8'h96] <= 32'h587c51b6 ;
    mem[8'h97] <= 32'h2dc21701 ;
    mem[8'h98] <= 32'hc189c8d2 ;
    mem[8'h99] <= 32'hb4378e65 ;
    mem[8'h9a] <= 32'h2af545bc ;
    mem[8'h9b] <= 32'h5f4b030b ;
    mem[8'h9c] <= 32'h13b1cfb9 ;
    mem[8'h9d] <= 32'h660f890e ;
    mem[8'h9e] <= 32'hf8cd42d7 ;
    mem[8'h9f] <= 32'h8d730460 ;
    mem[8'ha0] <= 32'hafdd962c ;
    mem[8'ha1] <= 32'hda63d09b ;
    mem[8'ha2] <= 32'h44a11b42 ;
    mem[8'ha3] <= 32'h311f5df5 ;
    mem[8'ha4] <= 32'h7de59147 ;
    mem[8'ha5] <= 32'h85bd7f0 ;
    mem[8'ha6] <= 32'h96991c29 ;
    mem[8'ha7] <= 32'he3275a9e ;
    mem[8'ha8] <= 32'hf6c854d ;
    mem[8'ha9] <= 32'h7ad2c3fa ;
    mem[8'haa] <= 32'he4100823 ;
    mem[8'hab] <= 32'h91ae4e94 ;
    mem[8'hac] <= 32'hdd548226 ;
    mem[8'had] <= 32'ha8eac491 ;
    mem[8'hae] <= 32'h36280f48 ;
    mem[8'haf] <= 32'h439649ff ;
    mem[8'hb0] <= 32'hea7ead59 ;
    mem[8'hb1] <= 32'h9fc0ebee ;
    mem[8'hb2] <= 32'h1022037 ;
    mem[8'hb3] <= 32'h74bc6680 ;
    mem[8'hb4] <= 32'h3846aa32 ;
    mem[8'hb5] <= 32'h4df8ec85 ;
    mem[8'hb6] <= 32'hd33a275c ;
    mem[8'hb7] <= 32'ha68461eb ;
    mem[8'hb8] <= 32'h4acfbe38 ;
    mem[8'hb9] <= 32'h3f71f88f ;
    mem[8'hba] <= 32'ha1b33356 ;
    mem[8'hbb] <= 32'hd40d75e1 ;
    mem[8'hbc] <= 32'h98f7b953 ;
    mem[8'hbd] <= 32'hed49ffe4 ;
    mem[8'hbe] <= 32'h738b343d ;
    mem[8'hbf] <= 32'h635728a ;
    mem[8'hc0] <= 32'h36d610a5 ;
    mem[8'hc1] <= 32'h43685612 ;
    mem[8'hc2] <= 32'hddaa9dcb ;
    mem[8'hc3] <= 32'ha814db7c ;
    mem[8'hc4] <= 32'he4ee17ce ;
    mem[8'hc5] <= 32'h91505179 ;
    mem[8'hc6] <= 32'hf929aa0 ;
    mem[8'hc7] <= 32'h7a2cdc17 ;
    mem[8'hc8] <= 32'h966703c4 ;
    mem[8'hc9] <= 32'he3d94573 ;
    mem[8'hca] <= 32'h7d1b8eaa ;
    mem[8'hcb] <= 32'h8a5c81d ;
    mem[8'hcc] <= 32'h445f04af ;
    mem[8'hcd] <= 32'h31e14218 ;
    mem[8'hce] <= 32'haf2389c1 ;
    mem[8'hcf] <= 32'hda9dcf76 ;
    mem[8'hd0] <= 32'h73752bd0 ;
    mem[8'hd1] <= 32'h6cb6d67 ;
    mem[8'hd2] <= 32'h9809a6be ;
    mem[8'hd3] <= 32'hedb7e009 ;
    mem[8'hd4] <= 32'ha14d2cbb ;
    mem[8'hd5] <= 32'hd4f36a0c ;
    mem[8'hd6] <= 32'h4a31a1d5 ;
    mem[8'hd7] <= 32'h3f8fe762 ;
    mem[8'hd8] <= 32'hd3c438b1 ;
    mem[8'hd9] <= 32'ha67a7e06 ;
    mem[8'hda] <= 32'h38b8b5df ;
    mem[8'hdb] <= 32'h4d06f368 ;
    mem[8'hdc] <= 32'h1fc3fda ;
    mem[8'hdd] <= 32'h7442796d ;
    mem[8'hde] <= 32'hea80b2b4 ;
    mem[8'hdf] <= 32'h9f3ef403 ;
    mem[8'he0] <= 32'hbd90664f ;
    mem[8'he1] <= 32'hc82e20f8 ;
    mem[8'he2] <= 32'h56eceb21 ;
    mem[8'he3] <= 32'h2352ad96 ;
    mem[8'he4] <= 32'h6fa86124 ;
    mem[8'he5] <= 32'h1a162793 ;
    mem[8'he6] <= 32'h84d4ec4a ;
    mem[8'he7] <= 32'hf16aaafd ;
    mem[8'he8] <= 32'h1d21752e ;
    mem[8'he9] <= 32'h689f3399 ;
    mem[8'hea] <= 32'hf65df840 ;
    mem[8'heb] <= 32'h83e3bef7 ;
    mem[8'hec] <= 32'hcf197245 ;
    mem[8'hed] <= 32'hbaa734f2 ;
    mem[8'hee] <= 32'h2465ff2b ;
    mem[8'hef] <= 32'h51dbb99c ;
    mem[8'hf0] <= 32'hf8335d3a ;
    mem[8'hf1] <= 32'h8d8d1b8d ;
    mem[8'hf2] <= 32'h134fd054 ;
    mem[8'hf3] <= 32'h66f196e3 ;
    mem[8'hf4] <= 32'h2a0b5a51 ;
    mem[8'hf5] <= 32'h5fb51ce6 ;
    mem[8'hf6] <= 32'hc177d73f ;
    mem[8'hf7] <= 32'hb4c99188 ;
    mem[8'hf8] <= 32'h58824e5b ;
    mem[8'hf9] <= 32'h2d3c08ec ;
    mem[8'hfa] <= 32'hb3fec335 ;
    mem[8'hfb] <= 32'hc6408582 ;
    mem[8'hfc] <= 32'h8aba4930 ;
    mem[8'hfd] <= 32'hff040f87 ;
    mem[8'hfe] <= 32'h61c6c45e ;
    mem[8'hff] <= 32'h147882e9 ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
