module crctab_ev19
(
input  wire         clk,
input  wire         rstn,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);
// ============================================================================
localparam  MEM_SIZE_BITS   = 8; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
// ============================================================================
wire [MEM_SIZE_BITS-1:0]    mem_addr;
wire [31:0]                 mem_data;
reg  [31:0]                 mem[0:MEM_SIZE];
initial begin
    mem[8'h0] <= 32'h0 ;
    mem[8'h1] <= 32'h34028fd6 ;
    mem[8'h2] <= 32'h68051fac ;
    mem[8'h3] <= 32'h5c07907a ;
    mem[8'h4] <= 32'hd00a3f58 ;
    mem[8'h5] <= 32'he408b08e ;
    mem[8'h6] <= 32'hb80f20f4 ;
    mem[8'h7] <= 32'h8c0daf22 ;
    mem[8'h8] <= 32'ha4d56307 ;
    mem[8'h9] <= 32'h90d7ecd1 ;
    mem[8'ha] <= 32'hccd07cab ;
    mem[8'hb] <= 32'hf8d2f37d ;
    mem[8'hc] <= 32'h74df5c5f ;
    mem[8'hd] <= 32'h40ddd389 ;
    mem[8'he] <= 32'h1cda43f3 ;
    mem[8'hf] <= 32'h28d8cc25 ;
    mem[8'h10] <= 32'h4d6bdbb9 ;
    mem[8'h11] <= 32'h7969546f ;
    mem[8'h12] <= 32'h256ec415 ;
    mem[8'h13] <= 32'h116c4bc3 ;
    mem[8'h14] <= 32'h9d61e4e1 ;
    mem[8'h15] <= 32'ha9636b37 ;
    mem[8'h16] <= 32'hf564fb4d ;
    mem[8'h17] <= 32'hc166749b ;
    mem[8'h18] <= 32'he9beb8be ;
    mem[8'h19] <= 32'hddbc3768 ;
    mem[8'h1a] <= 32'h81bba712 ;
    mem[8'h1b] <= 32'hb5b928c4 ;
    mem[8'h1c] <= 32'h39b487e6 ;
    mem[8'h1d] <= 32'hdb60830 ;
    mem[8'h1e] <= 32'h51b1984a ;
    mem[8'h1f] <= 32'h65b3179c ;
    mem[8'h20] <= 32'h9ad7b772 ;
    mem[8'h21] <= 32'haed538a4 ;
    mem[8'h22] <= 32'hf2d2a8de ;
    mem[8'h23] <= 32'hc6d02708 ;
    mem[8'h24] <= 32'h4add882a ;
    mem[8'h25] <= 32'h7edf07fc ;
    mem[8'h26] <= 32'h22d89786 ;
    mem[8'h27] <= 32'h16da1850 ;
    mem[8'h28] <= 32'h3e02d475 ;
    mem[8'h29] <= 32'ha005ba3 ;
    mem[8'h2a] <= 32'h5607cbd9 ;
    mem[8'h2b] <= 32'h6205440f ;
    mem[8'h2c] <= 32'hee08eb2d ;
    mem[8'h2d] <= 32'hda0a64fb ;
    mem[8'h2e] <= 32'h860df481 ;
    mem[8'h2f] <= 32'hb20f7b57 ;
    mem[8'h30] <= 32'hd7bc6ccb ;
    mem[8'h31] <= 32'he3bee31d ;
    mem[8'h32] <= 32'hbfb97367 ;
    mem[8'h33] <= 32'h8bbbfcb1 ;
    mem[8'h34] <= 32'h7b65393 ;
    mem[8'h35] <= 32'h33b4dc45 ;
    mem[8'h36] <= 32'h6fb34c3f ;
    mem[8'h37] <= 32'h5bb1c3e9 ;
    mem[8'h38] <= 32'h73690fcc ;
    mem[8'h39] <= 32'h476b801a ;
    mem[8'h3a] <= 32'h1b6c1060 ;
    mem[8'h3b] <= 32'h2f6e9fb6 ;
    mem[8'h3c] <= 32'ha3633094 ;
    mem[8'h3d] <= 32'h9761bf42 ;
    mem[8'h3e] <= 32'hcb662f38 ;
    mem[8'h3f] <= 32'hff64a0ee ;
    mem[8'h40] <= 32'h316e7353 ;
    mem[8'h41] <= 32'h56cfc85 ;
    mem[8'h42] <= 32'h596b6cff ;
    mem[8'h43] <= 32'h6d69e329 ;
    mem[8'h44] <= 32'he1644c0b ;
    mem[8'h45] <= 32'hd566c3dd ;
    mem[8'h46] <= 32'h896153a7 ;
    mem[8'h47] <= 32'hbd63dc71 ;
    mem[8'h48] <= 32'h95bb1054 ;
    mem[8'h49] <= 32'ha1b99f82 ;
    mem[8'h4a] <= 32'hfdbe0ff8 ;
    mem[8'h4b] <= 32'hc9bc802e ;
    mem[8'h4c] <= 32'h45b12f0c ;
    mem[8'h4d] <= 32'h71b3a0da ;
    mem[8'h4e] <= 32'h2db430a0 ;
    mem[8'h4f] <= 32'h19b6bf76 ;
    mem[8'h50] <= 32'h7c05a8ea ;
    mem[8'h51] <= 32'h4807273c ;
    mem[8'h52] <= 32'h1400b746 ;
    mem[8'h53] <= 32'h20023890 ;
    mem[8'h54] <= 32'hac0f97b2 ;
    mem[8'h55] <= 32'h980d1864 ;
    mem[8'h56] <= 32'hc40a881e ;
    mem[8'h57] <= 32'hf00807c8 ;
    mem[8'h58] <= 32'hd8d0cbed ;
    mem[8'h59] <= 32'hecd2443b ;
    mem[8'h5a] <= 32'hb0d5d441 ;
    mem[8'h5b] <= 32'h84d75b97 ;
    mem[8'h5c] <= 32'h8daf4b5 ;
    mem[8'h5d] <= 32'h3cd87b63 ;
    mem[8'h5e] <= 32'h60dfeb19 ;
    mem[8'h5f] <= 32'h54dd64cf ;
    mem[8'h60] <= 32'habb9c421 ;
    mem[8'h61] <= 32'h9fbb4bf7 ;
    mem[8'h62] <= 32'hc3bcdb8d ;
    mem[8'h63] <= 32'hf7be545b ;
    mem[8'h64] <= 32'h7bb3fb79 ;
    mem[8'h65] <= 32'h4fb174af ;
    mem[8'h66] <= 32'h13b6e4d5 ;
    mem[8'h67] <= 32'h27b46b03 ;
    mem[8'h68] <= 32'hf6ca726 ;
    mem[8'h69] <= 32'h3b6e28f0 ;
    mem[8'h6a] <= 32'h6769b88a ;
    mem[8'h6b] <= 32'h536b375c ;
    mem[8'h6c] <= 32'hdf66987e ;
    mem[8'h6d] <= 32'heb6417a8 ;
    mem[8'h6e] <= 32'hb76387d2 ;
    mem[8'h6f] <= 32'h83610804 ;
    mem[8'h70] <= 32'he6d21f98 ;
    mem[8'h71] <= 32'hd2d0904e ;
    mem[8'h72] <= 32'h8ed70034 ;
    mem[8'h73] <= 32'hbad58fe2 ;
    mem[8'h74] <= 32'h36d820c0 ;
    mem[8'h75] <= 32'h2daaf16 ;
    mem[8'h76] <= 32'h5edd3f6c ;
    mem[8'h77] <= 32'h6adfb0ba ;
    mem[8'h78] <= 32'h42077c9f ;
    mem[8'h79] <= 32'h7605f349 ;
    mem[8'h7a] <= 32'h2a026333 ;
    mem[8'h7b] <= 32'h1e00ece5 ;
    mem[8'h7c] <= 32'h920d43c7 ;
    mem[8'h7d] <= 32'ha60fcc11 ;
    mem[8'h7e] <= 32'hfa085c6b ;
    mem[8'h7f] <= 32'hce0ad3bd ;
    mem[8'h80] <= 32'h62dce6a6 ;
    mem[8'h81] <= 32'h56de6970 ;
    mem[8'h82] <= 32'had9f90a ;
    mem[8'h83] <= 32'h3edb76dc ;
    mem[8'h84] <= 32'hb2d6d9fe ;
    mem[8'h85] <= 32'h86d45628 ;
    mem[8'h86] <= 32'hdad3c652 ;
    mem[8'h87] <= 32'heed14984 ;
    mem[8'h88] <= 32'hc60985a1 ;
    mem[8'h89] <= 32'hf20b0a77 ;
    mem[8'h8a] <= 32'hae0c9a0d ;
    mem[8'h8b] <= 32'h9a0e15db ;
    mem[8'h8c] <= 32'h1603baf9 ;
    mem[8'h8d] <= 32'h2201352f ;
    mem[8'h8e] <= 32'h7e06a555 ;
    mem[8'h8f] <= 32'h4a042a83 ;
    mem[8'h90] <= 32'h2fb73d1f ;
    mem[8'h91] <= 32'h1bb5b2c9 ;
    mem[8'h92] <= 32'h47b222b3 ;
    mem[8'h93] <= 32'h73b0ad65 ;
    mem[8'h94] <= 32'hffbd0247 ;
    mem[8'h95] <= 32'hcbbf8d91 ;
    mem[8'h96] <= 32'h97b81deb ;
    mem[8'h97] <= 32'ha3ba923d ;
    mem[8'h98] <= 32'h8b625e18 ;
    mem[8'h99] <= 32'hbf60d1ce ;
    mem[8'h9a] <= 32'he36741b4 ;
    mem[8'h9b] <= 32'hd765ce62 ;
    mem[8'h9c] <= 32'h5b686140 ;
    mem[8'h9d] <= 32'h6f6aee96 ;
    mem[8'h9e] <= 32'h336d7eec ;
    mem[8'h9f] <= 32'h76ff13a ;
    mem[8'ha0] <= 32'hf80b51d4 ;
    mem[8'ha1] <= 32'hcc09de02 ;
    mem[8'ha2] <= 32'h900e4e78 ;
    mem[8'ha3] <= 32'ha40cc1ae ;
    mem[8'ha4] <= 32'h28016e8c ;
    mem[8'ha5] <= 32'h1c03e15a ;
    mem[8'ha6] <= 32'h40047120 ;
    mem[8'ha7] <= 32'h7406fef6 ;
    mem[8'ha8] <= 32'h5cde32d3 ;
    mem[8'ha9] <= 32'h68dcbd05 ;
    mem[8'haa] <= 32'h34db2d7f ;
    mem[8'hab] <= 32'hd9a2a9 ;
    mem[8'hac] <= 32'h8cd40d8b ;
    mem[8'had] <= 32'hb8d6825d ;
    mem[8'hae] <= 32'he4d11227 ;
    mem[8'haf] <= 32'hd0d39df1 ;
    mem[8'hb0] <= 32'hb5608a6d ;
    mem[8'hb1] <= 32'h816205bb ;
    mem[8'hb2] <= 32'hdd6595c1 ;
    mem[8'hb3] <= 32'he9671a17 ;
    mem[8'hb4] <= 32'h656ab535 ;
    mem[8'hb5] <= 32'h51683ae3 ;
    mem[8'hb6] <= 32'hd6faa99 ;
    mem[8'hb7] <= 32'h396d254f ;
    mem[8'hb8] <= 32'h11b5e96a ;
    mem[8'hb9] <= 32'h25b766bc ;
    mem[8'hba] <= 32'h79b0f6c6 ;
    mem[8'hbb] <= 32'h4db27910 ;
    mem[8'hbc] <= 32'hc1bfd632 ;
    mem[8'hbd] <= 32'hf5bd59e4 ;
    mem[8'hbe] <= 32'ha9bac99e ;
    mem[8'hbf] <= 32'h9db84648 ;
    mem[8'hc0] <= 32'h53b295f5 ;
    mem[8'hc1] <= 32'h67b01a23 ;
    mem[8'hc2] <= 32'h3bb78a59 ;
    mem[8'hc3] <= 32'hfb5058f ;
    mem[8'hc4] <= 32'h83b8aaad ;
    mem[8'hc5] <= 32'hb7ba257b ;
    mem[8'hc6] <= 32'hebbdb501 ;
    mem[8'hc7] <= 32'hdfbf3ad7 ;
    mem[8'hc8] <= 32'hf767f6f2 ;
    mem[8'hc9] <= 32'hc3657924 ;
    mem[8'hca] <= 32'h9f62e95e ;
    mem[8'hcb] <= 32'hab606688 ;
    mem[8'hcc] <= 32'h276dc9aa ;
    mem[8'hcd] <= 32'h136f467c ;
    mem[8'hce] <= 32'h4f68d606 ;
    mem[8'hcf] <= 32'h7b6a59d0 ;
    mem[8'hd0] <= 32'h1ed94e4c ;
    mem[8'hd1] <= 32'h2adbc19a ;
    mem[8'hd2] <= 32'h76dc51e0 ;
    mem[8'hd3] <= 32'h42dede36 ;
    mem[8'hd4] <= 32'hced37114 ;
    mem[8'hd5] <= 32'hfad1fec2 ;
    mem[8'hd6] <= 32'ha6d66eb8 ;
    mem[8'hd7] <= 32'h92d4e16e ;
    mem[8'hd8] <= 32'hba0c2d4b ;
    mem[8'hd9] <= 32'h8e0ea29d ;
    mem[8'hda] <= 32'hd20932e7 ;
    mem[8'hdb] <= 32'he60bbd31 ;
    mem[8'hdc] <= 32'h6a061213 ;
    mem[8'hdd] <= 32'h5e049dc5 ;
    mem[8'hde] <= 32'h2030dbf ;
    mem[8'hdf] <= 32'h36018269 ;
    mem[8'he0] <= 32'hc9652287 ;
    mem[8'he1] <= 32'hfd67ad51 ;
    mem[8'he2] <= 32'ha1603d2b ;
    mem[8'he3] <= 32'h9562b2fd ;
    mem[8'he4] <= 32'h196f1ddf ;
    mem[8'he5] <= 32'h2d6d9209 ;
    mem[8'he6] <= 32'h716a0273 ;
    mem[8'he7] <= 32'h45688da5 ;
    mem[8'he8] <= 32'h6db04180 ;
    mem[8'he9] <= 32'h59b2ce56 ;
    mem[8'hea] <= 32'h5b55e2c ;
    mem[8'heb] <= 32'h31b7d1fa ;
    mem[8'hec] <= 32'hbdba7ed8 ;
    mem[8'hed] <= 32'h89b8f10e ;
    mem[8'hee] <= 32'hd5bf6174 ;
    mem[8'hef] <= 32'he1bdeea2 ;
    mem[8'hf0] <= 32'h840ef93e ;
    mem[8'hf1] <= 32'hb00c76e8 ;
    mem[8'hf2] <= 32'hec0be692 ;
    mem[8'hf3] <= 32'hd8096944 ;
    mem[8'hf4] <= 32'h5404c666 ;
    mem[8'hf5] <= 32'h600649b0 ;
    mem[8'hf6] <= 32'h3c01d9ca ;
    mem[8'hf7] <= 32'h803561c ;
    mem[8'hf8] <= 32'h20db9a39 ;
    mem[8'hf9] <= 32'h14d915ef ;
    mem[8'hfa] <= 32'h48de8595 ;
    mem[8'hfb] <= 32'h7cdc0a43 ;
    mem[8'hfc] <= 32'hf0d1a561 ;
    mem[8'hfd] <= 32'hc4d32ab7 ;
    mem[8'hfe] <= 32'h98d4bacd ;
    mem[8'hff] <= 32'hacd6351b ;
end
assign mem_addr = addr[7:0];
// Output connectins
assign rdata    = mem_data;
assign mem_data = mem[mem_addr];
endmodule
